
library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

package CONV_PACK_overall is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_overall;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW01_add_25 is

   port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (29 downto 0);  CO : out std_logic);

end matrix_math_DW01_add_25;

architecture SYN_cla of matrix_math_DW01_add_25 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, SUM_14_port, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
      n54, n55, n56, n57, n58, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038 : std_logic;

begin
   SUM <= ( n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, A(13), A(12), A(11), A(10), A(9), 
      A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : INVX1 port map( A => n4, Y => n5);
   U3 : INVX1 port map( A => n58, Y => n6);
   U4 : INVX1 port map( A => n48, Y => n1);
   U5 : INVX2 port map( A => n45, Y => n48);
   U6 : INVX2 port map( A => n11, Y => n34);
   U7 : OR2X2 port map( A => A(18), B => B(18), Y => n33);
   U8 : XNOR2X1 port map( A => n28, B => n2, Y => SUM_20_port);
   U9 : NAND2X1 port map( A => n17, B => n22, Y => n2);
   U10 : AND2X2 port map( A => n52, B => n58, Y => SUM_14_port);
   U11 : INVX1 port map( A => n4, Y => n3);
   U12 : INVX2 port map( A => B(14), Y => n4);
   U13 : OR2X1 port map( A => n10, B => n3, Y => n52);
   U14 : NAND2X1 port map( A => n58, B => n7, Y => n8);
   U15 : NAND2X1 port map( A => n57, B => n6, Y => n9);
   U16 : NAND2X1 port map( A => n9, B => n8, Y => SUM_15_port);
   U17 : INVX1 port map( A => n57, Y => n7);
   U18 : BUFX2 port map( A => A(14), Y => n10);
   U19 : AND2X2 port map( A => n43, B => n1, Y => n11);
   U20 : AND2X2 port map( A => n11, B => n33, Y => n12);
   U21 : XNOR2X1 port map( A => n46, B => n47, Y => SUM_17_port);
   U22 : XNOR2X1 port map( A => n38, B => n39, Y => SUM_18_port);
   U23 : XNOR2X1 port map( A => n30, B => n31, Y => SUM_19_port);
   U24 : NAND2X1 port map( A => n49, B => n50, Y => n25);
   U25 : NAND2X1 port map( A => n56, B => n50, Y => n54);
   U26 : XOR2X1 port map( A => n14, B => n15, Y => SUM_21_port);
   U27 : XOR2X1 port map( A => B(21), B => A(21), Y => n15);
   U28 : NAND2X1 port map( A => n16, B => n17, Y => n14);
   U29 : OAI21X1 port map( A => n18, B => n19, C => n20, Y => n16);
   U30 : AND2X2 port map( A => n21, B => n22, Y => n20);
   U31 : NAND2X1 port map( A => n23, B => n24, Y => n19);
   U32 : NAND2X1 port map( A => n12, B => n25, Y => n24);
   U33 : NAND2X1 port map( A => n26, B => n27, Y => n18);
   U34 : OR2X2 port map( A => A(20), B => B(20), Y => n22);
   U35 : NAND2X1 port map( A => B(20), B => A(20), Y => n17);
   U36 : NAND2X1 port map( A => n29, B => n27, Y => n28);
   U37 : NAND2X1 port map( A => n21, B => n30, Y => n29);
   U38 : NAND2X1 port map( A => n27, B => n21, Y => n31);
   U39 : OR2X2 port map( A => A(19), B => B(19), Y => n21);
   U40 : NAND2X1 port map( A => B(19), B => A(19), Y => n27);
   U41 : NAND3X1 port map( A => n23, B => n26, C => n32, Y => n30);
   U42 : NAND2X1 port map( A => n25, B => n12, Y => n32);
   U43 : NAND2X1 port map( A => n35, B => n33, Y => n23);
   U44 : NAND2X1 port map( A => n36, B => n37, Y => n35);
   U45 : NAND2X1 port map( A => n26, B => n33, Y => n39);
   U46 : NAND2X1 port map( A => A(18), B => B(18), Y => n26);
   U47 : OAI21X1 port map( A => n40, B => n34, C => n41, Y => n38);
   U48 : AND2X2 port map( A => n36, B => n37, Y => n41);
   U49 : NAND2X1 port map( A => n43, B => n42, Y => n36);
   U50 : INVX2 port map( A => n44, Y => n42);
   U51 : NAND2X1 port map( A => n43, B => n37, Y => n47);
   U52 : OR2X2 port map( A => A(17), B => B(17), Y => n43);
   U53 : NAND2X1 port map( A => A(17), B => B(17), Y => n37);
   U54 : OAI21X1 port map( A => n40, B => n48, C => n44, Y => n46);
   U55 : INVX2 port map( A => n25, Y => n40);
   U56 : NAND2X1 port map( A => n51, B => n53, Y => n49);
   U57 : AND2X2 port map( A => B(14), B => A(14), Y => n53);
   U58 : XNOR2X1 port map( A => n54, B => n55, Y => SUM_16_port);
   U59 : NAND2X1 port map( A => n45, B => n44, Y => n55);
   U60 : NAND2X1 port map( A => A(16), B => B(16), Y => n44);
   U61 : OR2X2 port map( A => B(16), B => A(16), Y => n45);
   U62 : NAND2X1 port map( A => n51, B => n53, Y => n56);
   U63 : NAND2X1 port map( A => n51, B => n50, Y => n57);
   U64 : NAND2X1 port map( A => A(15), B => B(15), Y => n50);
   U65 : OR2X2 port map( A => A(15), B => B(15), Y => n51);
   U66 : NAND2X1 port map( A => n5, B => n10, Y => n58);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW01_add_24 is

   port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (29 downto 0);  CO : out std_logic);

end matrix_math_DW01_add_24;

architecture SYN_cla of matrix_math_DW01_add_24 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, SUM_14_port, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078 : std_logic;

begin
   SUM <= ( n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, A(13), A(12), A(11), A(10), A(9), 
      A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2X2 port map( A => A(17), B => B(17), Y => n1);
   U3 : BUFX2 port map( A => A(14), Y => n2);
   U4 : BUFX2 port map( A => B(14), Y => n3);
   U5 : OR2X1 port map( A => n2, B => n3, Y => n43);
   U6 : XOR2X1 port map( A => n4, B => n24, Y => SUM_19_port);
   U7 : INVX1 port map( A => n22, Y => n4);
   U8 : OR2X2 port map( A => A(15), B => B(15), Y => n8);
   U9 : XNOR2X1 port map( A => n38, B => n5, Y => SUM_17_port);
   U10 : NAND2X1 port map( A => n1, B => n36, Y => n5);
   U11 : NOR2X1 port map( A => A(17), B => B(17), Y => n6);
   U12 : AND2X2 port map( A => n10, B => n1, Y => n7);
   U13 : INVX1 port map( A => n39, Y => n10);
   U14 : OR2X1 port map( A => A(15), B => B(15), Y => n42);
   U15 : XNOR2X1 port map( A => n9, B => n44, Y => SUM_16_port);
   U16 : NAND2X1 port map( A => n45, B => n41, Y => n9);
   U17 : INVX1 port map( A => n37, Y => n39);
   U18 : AND2X2 port map( A => A(14), B => B(14), Y => n46);
   U19 : XOR2X1 port map( A => n14, B => n11, Y => SUM_21_port);
   U20 : XNOR2X1 port map( A => B(21), B => A(21), Y => n11);
   U21 : XNOR2X1 port map( A => n32, B => n33, Y => SUM_18_port);
   U22 : XOR2X1 port map( A => n48, B => n47, Y => SUM_15_port);
   U23 : AND2X2 port map( A => n40, B => n41, Y => n12);
   U24 : AND2X2 port map( A => n43, B => n48, Y => SUM_14_port);
   U25 : AOI21X1 port map( A => n20, B => n15, C => n16, Y => n14);
   U26 : INVX2 port map( A => n17, Y => n16);
   U27 : XNOR2X1 port map( A => n21, B => n20, Y => SUM_20_port);
   U28 : NAND2X1 port map( A => n15, B => n17, Y => n21);
   U29 : NAND2X1 port map( A => B(20), B => A(20), Y => n17);
   U30 : OR2X2 port map( A => A(20), B => B(20), Y => n15);
   U31 : NAND2X1 port map( A => n19, B => n18, Y => n20);
   U32 : NAND2X1 port map( A => n22, B => n23, Y => n19);
   U33 : NAND2X1 port map( A => n23, B => n18, Y => n24);
   U34 : NAND2X1 port map( A => A(19), B => B(19), Y => n18);
   U35 : OR2X2 port map( A => A(19), B => B(19), Y => n23);
   U36 : OAI21X1 port map( A => n12, B => n25, C => n26, Y => n22);
   U37 : AOI21X1 port map( A => n28, B => n27, C => n29, Y => n26);
   U38 : INVX2 port map( A => n30, Y => n29);
   U39 : NAND2X1 port map( A => n28, B => n7, Y => n25);
   U40 : NAND2X1 port map( A => n30, B => n28, Y => n33);
   U41 : OR2X2 port map( A => A(18), B => B(18), Y => n28);
   U42 : NAND2X1 port map( A => B(18), B => A(18), Y => n30);
   U43 : OAI21X1 port map( A => n12, B => n31, C => n34, Y => n32);
   U44 : INVX2 port map( A => n27, Y => n34);
   U45 : OAI21X1 port map( A => n6, B => n35, C => n36, Y => n27);
   U46 : NAND2X1 port map( A => n10, B => n1, Y => n31);
   U47 : NAND2X1 port map( A => A(17), B => B(17), Y => n36);
   U48 : OAI21X1 port map( A => n39, B => n12, C => n35, Y => n38);
   U49 : NAND2X1 port map( A => n8, B => n46, Y => n40);
   U50 : NAND2X1 port map( A => n35, B => n37, Y => n44);
   U51 : NAND2X1 port map( A => A(16), B => B(16), Y => n35);
   U52 : OR2X2 port map( A => A(16), B => B(16), Y => n37);
   U53 : NAND2X1 port map( A => n42, B => n46, Y => n45);
   U54 : NAND2X1 port map( A => n41, B => n8, Y => n47);
   U55 : NAND2X1 port map( A => A(15), B => B(15), Y => n41);
   U56 : NAND2X1 port map( A => n3, B => n2, Y => n48);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW01_add_23 is

   port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (29 downto 0);  CO : out std_logic);

end matrix_math_DW01_add_23;

architecture SYN_cla of matrix_math_DW01_add_23 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, SUM_14_port, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
      n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n_1111, n_1112, 
      n_1113, n_1114, n_1115, n_1116, n_1117, n_1118 : std_logic;

begin
   SUM <= ( n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, A(13), A(12), A(11), A(10), A(9), 
      A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : AND2X2 port map( A => n20, B => n29, Y => n2);
   U3 : OR2X1 port map( A => B(16), B => A(16), Y => n1);
   U4 : OR2X1 port map( A => A(16), B => B(16), Y => n54);
   U5 : AND2X1 port map( A => n29, B => n30, Y => n28);
   U6 : INVX2 port map( A => n44, Y => n34);
   U7 : INVX1 port map( A => n31, Y => n26);
   U8 : NAND2X1 port map( A => n3, B => n2, Y => n4);
   U9 : NAND2X1 port map( A => n4, B => n35, Y => n32);
   U10 : INVX1 port map( A => n34, Y => n3);
   U11 : INVX1 port map( A => n27, Y => n5);
   U12 : INVX1 port map( A => n5, Y => n6);
   U13 : INVX1 port map( A => A(14), Y => n7);
   U14 : INVX1 port map( A => n7, Y => n8);
   U15 : OR2X1 port map( A => n16, B => n13, Y => n60);
   U16 : XNOR2X1 port map( A => n50, B => n9, Y => SUM_18_port);
   U17 : NAND2X1 port map( A => n40, B => n45, Y => n9);
   U18 : INVX1 port map( A => A(19), Y => n10);
   U19 : INVX1 port map( A => n10, Y => n11);
   U20 : OR2X2 port map( A => A(15), B => B(15), Y => n12);
   U21 : OR2X1 port map( A => A(15), B => B(15), Y => n59);
   U22 : INVX1 port map( A => n41, Y => n36);
   U23 : BUFX2 port map( A => B(14), Y => n13);
   U24 : BUFX2 port map( A => n1, Y => n14);
   U25 : AND2X2 port map( A => n53, B => n1, Y => n15);
   U26 : INVX1 port map( A => n15, Y => n46);
   U27 : BUFX2 port map( A => A(14), Y => n16);
   U28 : XNOR2X1 port map( A => n62, B => n17, Y => SUM_16_port);
   U29 : NAND2X1 port map( A => n56, B => n54, Y => n17);
   U30 : XOR2X1 port map( A => n64, B => n18, Y => SUM_15_port);
   U31 : NAND2X1 port map( A => n58, B => n12, Y => n18);
   U32 : XNOR2X1 port map( A => n55, B => n19, Y => SUM_17_port);
   U33 : AND2X2 port map( A => n49, B => n53, Y => n19);
   U34 : AND2X2 port map( A => n15, B => n45, Y => n20);
   U35 : XNOR2X1 port map( A => n27, B => n42, Y => SUM_19_port);
   U36 : AND2X2 port map( A => n64, B => n60, Y => SUM_14_port);
   U37 : NAND2X1 port map( A => n57, B => n58, Y => n44);
   U38 : NAND2X1 port map( A => n58, B => n63, Y => n62);
   U39 : XOR2X1 port map( A => n22, B => n23, Y => SUM_21_port);
   U40 : XOR2X1 port map( A => B(21), B => A(21), Y => n23);
   U41 : NAND2X1 port map( A => n24, B => n25, Y => n22);
   U42 : OAI21X1 port map( A => n26, B => n6, C => n28, Y => n25);
   U43 : XNOR2X1 port map( A => n32, B => n33, Y => SUM_20_port);
   U44 : NAND2X1 port map( A => n30, B => n24, Y => n33);
   U45 : NAND2X1 port map( A => B(20), B => A(20), Y => n24);
   U46 : OR2X2 port map( A => A(20), B => B(20), Y => n30);
   U47 : AOI21X1 port map( A => n36, B => n29, C => n37, Y => n35);
   U48 : NAND2X1 port map( A => n31, B => n38, Y => n37);
   U49 : NAND2X1 port map( A => n39, B => n29, Y => n38);
   U50 : INVX2 port map( A => n40, Y => n39);
   U51 : NAND2X1 port map( A => n31, B => n29, Y => n42);
   U52 : OR2X2 port map( A => A(19), B => B(19), Y => n29);
   U53 : NAND2X1 port map( A => n11, B => B(19), Y => n31);
   U54 : NAND3X1 port map( A => n41, B => n40, C => n43, Y => n27);
   U55 : NAND2X1 port map( A => n44, B => n20, Y => n43);
   U56 : NAND2X1 port map( A => n47, B => n45, Y => n41);
   U57 : NAND2X1 port map( A => n48, B => n49, Y => n47);
   U58 : OR2X2 port map( A => A(18), B => B(18), Y => n45);
   U59 : NAND2X1 port map( A => B(18), B => A(18), Y => n40);
   U60 : OAI21X1 port map( A => n34, B => n46, C => n51, Y => n50);
   U61 : AND2X2 port map( A => n48, B => n49, Y => n51);
   U62 : NAND2X1 port map( A => n53, B => n52, Y => n48);
   U63 : OR2X2 port map( A => A(17), B => B(17), Y => n53);
   U64 : NAND2X1 port map( A => B(17), B => A(17), Y => n49);
   U65 : AOI21X1 port map( A => n44, B => n14, C => n52, Y => n55);
   U66 : INVX2 port map( A => n56, Y => n52);
   U67 : NAND2X1 port map( A => n12, B => n61, Y => n57);
   U68 : AND2X2 port map( A => A(14), B => B(14), Y => n61);
   U69 : NAND2X1 port map( A => A(16), B => B(16), Y => n56);
   U70 : NAND2X1 port map( A => n59, B => n61, Y => n63);
   U71 : NAND2X1 port map( A => A(15), B => B(15), Y => n58);
   U72 : NAND2X1 port map( A => n8, B => n13, Y => n64);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW01_add_18 is

   port( A, B : in std_logic_vector (23 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (23 downto 0);  CO : out std_logic);

end matrix_math_DW01_add_18;

architecture SYN_cla of matrix_math_DW01_add_18 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132 : std_logic;

begin
   
   U2 : INVX1 port map( A => A(19), Y => n1);
   U3 : INVX1 port map( A => n1, Y => n2);
   U4 : INVX1 port map( A => n22, Y => n3);
   U5 : BUFX2 port map( A => n61, Y => n4);
   U6 : INVX1 port map( A => n56, Y => n13);
   U7 : INVX1 port map( A => n21, Y => n5);
   U8 : INVX2 port map( A => A(18), Y => n21);
   U9 : INVX1 port map( A => n47, Y => n6);
   U10 : INVX1 port map( A => n47, Y => n33);
   U11 : AND2X1 port map( A => B(21), B => n8, Y => n28);
   U12 : INVX1 port map( A => A(21), Y => n7);
   U13 : INVX1 port map( A => n7, Y => n8);
   U14 : OR2X2 port map( A => A(19), B => B(19), Y => n9);
   U15 : OR2X1 port map( A => A(19), B => B(19), Y => n29);
   U16 : AND2X1 port map( A => B(19), B => A(19), Y => n64);
   U17 : INVX1 port map( A => A(20), Y => n10);
   U18 : INVX1 port map( A => A(20), Y => n23);
   U19 : INVX1 port map( A => n48, Y => n11);
   U20 : NAND2X1 port map( A => n23, B => n24, Y => n12);
   U21 : INVX2 port map( A => B(20), Y => n24);
   U22 : XOR2X1 port map( A => n13, B => n57, Y => SUM(21));
   U23 : INVX2 port map( A => n14, Y => n44);
   U24 : NAND3X1 port map( A => n29, B => n58, C => n59, Y => n14);
   U25 : INVX2 port map( A => n75, Y => n19);
   U26 : INVX2 port map( A => n25, Y => n26);
   U27 : NAND2X1 port map( A => B(7), B => A(7), Y => n15);
   U28 : AND2X2 port map( A => B(3), B => A(3), Y => n16);
   U29 : NOR2X1 port map( A => A(3), B => B(3), Y => n17);
   U30 : NOR2X1 port map( A => A(1), B => B(1), Y => n18);
   U31 : XOR2X1 port map( A => n76, B => n19, Y => SUM(18));
   U32 : XNOR2X1 port map( A => n65, B => n66, Y => SUM(20));
   U33 : XOR2X1 port map( A => n54, B => n55, Y => SUM(22));
   U34 : INVX1 port map( A => n23, Y => n20);
   U35 : NAND2X1 port map( A => n22, B => n21, Y => n73);
   U36 : INVX1 port map( A => B(18), Y => n22);
   U37 : NAND2X1 port map( A => n24, B => n10, Y => n58);
   U38 : INVX1 port map( A => B(20), Y => n25);
   U39 : BUFX2 port map( A => n62, Y => n27);
   U40 : AND2X1 port map( A => B(17), B => A(17), Y => n74);
   U41 : BUFX2 port map( A => n5, Y => n30);
   U42 : BUFX2 port map( A => n63, Y => n31);
   U43 : BUFX2 port map( A => n3, Y => n32);
   U44 : XNOR2X1 port map( A => n41, B => n34, Y => SUM(23));
   U45 : XNOR2X1 port map( A => A(23), B => B(23), Y => n34);
   U46 : INVX1 port map( A => n48, Y => n35);
   U47 : NOR2X1 port map( A => A(21), B => B(21), Y => n36);
   U48 : INVX1 port map( A => n36, Y => n49);
   U49 : AND2X1 port map( A => n72, B => n77, Y => n37);
   U50 : AND2X2 port map( A => B(14), B => A(14), Y => n38);
   U51 : AND2X2 port map( A => B(12), B => A(12), Y => n39);
   U52 : AND2X2 port map( A => B(10), B => A(10), Y => n40);
   U53 : AND2X1 port map( A => n63, B => n62, Y => n60);
   U54 : NAND2X1 port map( A => n42, B => n43, Y => n41);
   U55 : OAI21X1 port map( A => n44, B => n45, C => n46, Y => n43);
   U56 : AOI21X1 port map( A => n47, B => n48, C => n36, Y => n46);
   U57 : INVX2 port map( A => B(22), Y => n48);
   U58 : INVX2 port map( A => A(22), Y => n47);
   U59 : NAND3X1 port map( A => n50, B => n51, C => n52, Y => n45);
   U60 : NAND2X1 port map( A => A(21), B => B(21), Y => n51);
   U61 : OAI21X1 port map( A => n33, B => n35, C => n42, Y => n55);
   U62 : NAND2X1 port map( A => n6, B => n11, Y => n42);
   U63 : AOI21X1 port map( A => n56, B => n49, C => n28, Y => n54);
   U64 : NAND2X1 port map( A => n51, B => n49, Y => n57);
   U65 : NAND3X1 port map( A => n50, B => n52, C => n53, Y => n56);
   U66 : NAND3X1 port map( A => n9, B => n12, C => n59, Y => n53);
   U67 : NAND2X1 port map( A => n60, B => n61, Y => n59);
   U68 : OAI21X1 port map( A => A(20), B => B(20), C => n64, Y => n50);
   U69 : OAI21X1 port map( A => n20, B => n26, C => n52, Y => n66);
   U70 : NAND2X1 port map( A => A(20), B => B(20), Y => n52);
   U71 : NAND2X1 port map( A => n67, B => n68, Y => n65);
   U72 : NAND2X1 port map( A => n9, B => n69, Y => n68);
   U73 : XNOR2X1 port map( A => n70, B => n69, Y => SUM(19));
   U74 : NAND2X1 port map( A => n67, B => n9, Y => n70);
   U75 : NAND2X1 port map( A => B(19), B => n2, Y => n67);
   U76 : NAND3X1 port map( A => n31, B => n27, C => n4, Y => n69);
   U77 : NAND3X1 port map( A => n71, B => n72, C => n73, Y => n61);
   U78 : OAI21X1 port map( A => B(18), B => A(18), C => n74, Y => n62);
   U79 : OAI21X1 port map( A => n30, B => n32, C => n31, Y => n76);
   U80 : NAND2X1 port map( A => A(18), B => B(18), Y => n63);
   U81 : NAND2X1 port map( A => n77, B => n78, Y => n75);
   U82 : NAND2X1 port map( A => n71, B => n72, Y => n78);
   U83 : NAND2X1 port map( A => n79, B => n80, Y => n71);
   U84 : OAI21X1 port map( A => A(16), B => B(16), C => n81, Y => n80);
   U85 : NAND2X1 port map( A => A(16), B => B(16), Y => n79);
   U86 : XOR2X1 port map( A => n82, B => n37, Y => SUM(17));
   U87 : NAND2X1 port map( A => B(17), B => A(17), Y => n77);
   U88 : OR2X2 port map( A => B(17), B => A(17), Y => n72);
   U89 : NAND2X1 port map( A => n83, B => n84, Y => n82);
   U90 : OAI21X1 port map( A => B(16), B => A(16), C => n81, Y => n84);
   U91 : XNOR2X1 port map( A => n81, B => n85, Y => SUM(16));
   U92 : OAI21X1 port map( A => A(16), B => B(16), C => n83, Y => n85);
   U93 : NAND2X1 port map( A => B(16), B => A(16), Y => n83);
   U94 : OAI22X1 port map( A => n86, B => n87, C => n88, D => n89, Y => n81);
   U95 : OAI21X1 port map( A => n38, B => n90, C => n91, Y => n89);
   U96 : OR2X2 port map( A => A(14), B => B(14), Y => n91);
   U97 : OAI21X1 port map( A => n92, B => n93, C => n94, Y => n90);
   U98 : NAND2X1 port map( A => B(13), B => A(13), Y => n94);
   U99 : OAI21X1 port map( A => n39, B => n95, C => n96, Y => n93);
   U100 : OR2X2 port map( A => A(12), B => B(12), Y => n96);
   U101 : OAI22X1 port map( A => n97, B => n98, C => n99, D => n100, Y => n95);
   U102 : OAI21X1 port map( A => n101, B => n40, C => n102, Y => n100);
   U103 : OR2X2 port map( A => A(10), B => B(10), Y => n102);
   U104 : NAND3X1 port map( A => n103, B => n104, C => n105, Y => n101);
   U105 : NAND2X1 port map( A => B(9), B => A(9), Y => n105);
   U106 : NAND3X1 port map( A => n106, B => n107, C => n108, Y => n104);
   U107 : AOI22X1 port map( A => n109, B => n110, C => n111, D => n112, Y => 
                           n107);
   U108 : INVX2 port map( A => A(8), Y => n112);
   U109 : INVX2 port map( A => B(8), Y => n111);
   U110 : INVX2 port map( A => A(7), Y => n110);
   U111 : INVX2 port map( A => B(7), Y => n109);
   U112 : NAND3X1 port map( A => n113, B => n114, C => n15, Y => n106);
   U113 : OAI21X1 port map( A => n117, B => n16, C => n115, Y => n114);
   U114 : INVX2 port map( A => n118, Y => n115);
   U115 : NAND3X1 port map( A => n119, B => n120, C => n121, Y => n118);
   U116 : OR2X2 port map( A => A(4), B => B(4), Y => n119);
   U117 : AOI21X1 port map( A => n122, B => n123, C => n17, Y => n117);
   U118 : NAND2X1 port map( A => n124, B => n116, Y => n123);
   U119 : OR2X2 port map( A => A(2), B => B(2), Y => n116);
   U120 : OAI22X1 port map( A => n125, B => n126, C => n18, D => n127, Y => 
                           n124);
   U121 : NAND2X1 port map( A => A(0), B => B(0), Y => n127);
   U122 : INVX2 port map( A => B(1), Y => n126);
   U123 : INVX2 port map( A => A(1), Y => n125);
   U124 : NAND2X1 port map( A => B(2), B => A(2), Y => n122);
   U125 : AOI22X1 port map( A => B(6), B => A(6), C => n128, D => n121, Y => 
                           n113);
   U126 : OR2X2 port map( A => A(6), B => B(6), Y => n121);
   U127 : AOI21X1 port map( A => n129, B => n130, C => n131, Y => n128);
   U128 : INVX2 port map( A => n120, Y => n131);
   U129 : OR2X2 port map( A => A(5), B => B(5), Y => n120);
   U130 : NAND2X1 port map( A => B(5), B => A(5), Y => n130);
   U131 : NAND2X1 port map( A => B(4), B => A(4), Y => n129);
   U132 : NAND2X1 port map( A => n132, B => n108, Y => n103);
   U133 : OR2X2 port map( A => A(9), B => B(9), Y => n108);
   U134 : AND2X2 port map( A => A(8), B => B(8), Y => n132);
   U135 : NOR2X1 port map( A => A(11), B => B(11), Y => n99);
   U136 : INVX2 port map( A => B(11), Y => n98);
   U137 : INVX2 port map( A => A(11), Y => n97);
   U138 : NOR2X1 port map( A => A(13), B => B(13), Y => n92);
   U139 : NOR2X1 port map( A => A(15), B => B(15), Y => n88);
   U140 : INVX2 port map( A => B(15), Y => n87);
   U141 : INVX2 port map( A => A(15), Y => n86);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW01_add_13 is

   port( A, B : in std_logic_vector (23 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (23 downto 0);  CO : out std_logic);

end matrix_math_DW01_add_13;

architecture SYN_cla of matrix_math_DW01_add_13 is

   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160 : std_logic;

begin
   
   U2 : NAND3X1 port map( A => n74, B => n73, C => n72, Y => n1);
   U3 : OR2X1 port map( A => A(22), B => B(22), Y => n66);
   U4 : AND2X2 port map( A => A(22), B => B(22), Y => n6);
   U5 : XNOR2X1 port map( A => n13, B => n2, Y => SUM(21));
   U6 : NAND2X1 port map( A => n79, B => n72, Y => n2);
   U7 : NAND2X1 port map( A => n3, B => n4, Y => n5);
   U8 : NAND2X1 port map( A => n5, B => n101, Y => n100);
   U9 : INVX1 port map( A => n19, Y => n3);
   U10 : INVX2 port map( A => n98, Y => n4);
   U11 : AND2X2 port map( A => n87, B => n86, Y => SUM(0));
   U12 : XNOR2X1 port map( A => A(22), B => B(22), Y => n67);
   U13 : AND2X1 port map( A => n103, B => n10, Y => n101);
   U14 : NOR2X1 port map( A => B(17), B => A(17), Y => n8);
   U15 : INVX2 port map( A => n26, Y => n27);
   U16 : OAI21X1 port map( A => n69, B => n70, C => n71, Y => n9);
   U17 : OR2X2 port map( A => B(17), B => A(17), Y => n10);
   U18 : BUFX2 port map( A => A(18), Y => n11);
   U19 : XOR2X1 port map( A => n64, B => n12, Y => SUM(23));
   U20 : XNOR2X1 port map( A => B(23), B => A(23), Y => n12);
   U21 : NAND2X1 port map( A => n71, B => n74, Y => n13);
   U22 : XOR2X1 port map( A => n99, B => n14, Y => SUM(18));
   U23 : AND2X2 port map( A => n94, B => n93, Y => n14);
   U24 : XOR2X1 port map( A => n67, B => n9, Y => SUM(22));
   U25 : NOR2X1 port map( A => n15, B => n8, Y => n90);
   U26 : INVX1 port map( A => n15, Y => n94);
   U27 : NOR2X1 port map( A => A(18), B => B(18), Y => n15);
   U28 : AND2X2 port map( A => B(16), B => A(16), Y => n19);
   U29 : INVX1 port map( A => n137, Y => n147);
   U30 : INVX1 port map( A => n42, Y => n41);
   U31 : XOR2X1 port map( A => n83, B => n84, Y => SUM(20));
   U32 : XOR2X1 port map( A => n27, B => n88, Y => SUM(19));
   U33 : XOR2X1 port map( A => n102, B => n17, Y => SUM(17));
   U34 : NAND2X1 port map( A => n10, B => n92, Y => n17);
   U35 : XNOR2X1 port map( A => n124, B => n125, Y => SUM(15));
   U36 : XNOR2X1 port map( A => n127, B => n18, Y => SUM(14));
   U37 : NAND2X1 port map( A => n107, B => n112, Y => n18);
   U38 : XOR2X1 port map( A => n104, B => n98, Y => SUM(16));
   U39 : XOR2X1 port map( A => n133, B => n20, Y => SUM(12));
   U40 : NAND2X1 port map( A => n122, B => n117, Y => n20);
   U41 : XOR2X1 port map( A => n144, B => n145, Y => SUM(11));
   U42 : NOR2X1 port map( A => n142, B => n143, Y => n21);
   U43 : XNOR2X1 port map( A => n146, B => n22, Y => SUM(10));
   U44 : NAND2X1 port map( A => n141, B => n137, Y => n22);
   U45 : XOR2X1 port map( A => n28, B => n23, Y => SUM(9));
   U46 : NAND2X1 port map( A => n29, B => n30, Y => n23);
   U47 : XNOR2X1 port map( A => n39, B => n24, Y => SUM(6));
   U48 : NAND2X1 port map( A => n40, B => n42, Y => n24);
   U49 : XNOR2X1 port map( A => n31, B => n32, Y => SUM(8));
   U50 : XOR2X1 port map( A => n35, B => n36, Y => SUM(7));
   U51 : XNOR2X1 port map( A => n45, B => n25, Y => SUM(5));
   U52 : NAND2X1 port map( A => n46, B => n44, Y => n25);
   U53 : INVX2 port map( A => n86, Y => n62);
   U54 : NAND2X1 port map( A => n115, B => n116, Y => n114);
   U55 : INVX2 port map( A => n81, Y => n26);
   U56 : NAND2X1 port map( A => n33, B => n34, Y => n32);
   U57 : NAND2X1 port map( A => n37, B => n38, Y => n36);
   U58 : AOI21X1 port map( A => n39, B => n40, C => n41, Y => n35);
   U59 : NAND2X1 port map( A => n43, B => n44, Y => n39);
   U60 : NAND2X1 port map( A => n45, B => n46, Y => n43);
   U61 : OAI21X1 port map( A => n119, B => n47, C => n48, Y => n45);
   U62 : INVX2 port map( A => n49, Y => n47);
   U63 : XNOR2X1 port map( A => n50, B => n155, Y => SUM(4));
   U64 : NAND2X1 port map( A => n48, B => n49, Y => n50);
   U65 : XNOR2X1 port map( A => n51, B => n52, Y => SUM(3));
   U66 : AND2X2 port map( A => n53, B => n54, Y => n52);
   U67 : AOI21X1 port map( A => n55, B => n56, C => n57, Y => n51);
   U68 : INVX2 port map( A => n58, Y => n57);
   U69 : XNOR2X1 port map( A => n59, B => n60, Y => SUM(2));
   U70 : AND2X2 port map( A => n56, B => n58, Y => n60);
   U71 : INVX2 port map( A => n55, Y => n59);
   U72 : OAI21X1 port map( A => n160, B => n86, C => n61, Y => n55);
   U73 : AOI21X1 port map( A => n66, B => n65, C => n6, Y => n64);
   U74 : INVX2 port map( A => n68, Y => n65);
   U75 : OAI21X1 port map( A => n69, B => n1, C => n71, Y => n68);
   U76 : NAND3X1 port map( A => n74, B => n73, C => n72, Y => n70);
   U77 : NAND2X1 port map( A => n76, B => n75, Y => n73);
   U78 : INVX2 port map( A => n77, Y => n69);
   U79 : NAND3X1 port map( A => n78, B => n76, C => n26, Y => n77);
   U80 : NAND2X1 port map( A => B(21), B => A(21), Y => n74);
   U81 : OR2X2 port map( A => A(21), B => B(21), Y => n71);
   U82 : NAND3X1 port map( A => n78, B => n76, C => n80, Y => n79);
   U83 : NAND2X1 port map( A => n82, B => n81, Y => n80);
   U84 : NAND2X1 port map( A => n72, B => n76, Y => n84);
   U85 : OR2X2 port map( A => A(20), B => B(20), Y => n76);
   U86 : NAND2X1 port map( A => B(20), B => A(20), Y => n72);
   U87 : AOI21X1 port map( A => n26, B => n78, C => n75, Y => n83);
   U88 : INVX2 port map( A => n82, Y => n75);
   U89 : XNOR2X1 port map( A => n85, B => n62, Y => SUM(1));
   U90 : NAND2X1 port map( A => n63, B => n61, Y => n85);
   U91 : AOI21X1 port map( A => n89, B => n90, C => n91, Y => n81);
   U92 : OAI21X1 port map( A => n15, B => n92, C => n93, Y => n91);
   U93 : AOI21X1 port map( A => n95, B => n96, C => n97, Y => n89);
   U94 : NOR2X1 port map( A => B(16), B => A(16), Y => n97);
   U95 : INVX2 port map( A => n98, Y => n96);
   U96 : NAND2X1 port map( A => B(16), B => A(16), Y => n95);
   U97 : NAND2X1 port map( A => n82, B => n78, Y => n88);
   U98 : OR2X2 port map( A => B(19), B => A(19), Y => n78);
   U99 : NAND2X1 port map( A => B(19), B => A(19), Y => n82);
   U100 : NAND2X1 port map( A => n11, B => B(18), Y => n93);
   U101 : NAND2X1 port map( A => n92, B => n100, Y => n99);
   U102 : NAND2X1 port map( A => B(17), B => A(17), Y => n92);
   U103 : AOI21X1 port map( A => n98, B => n103, C => n19, Y => n102);
   U104 : OR2X2 port map( A => A(16), B => B(16), Y => n103);
   U105 : NAND2X1 port map( A => n105, B => n106, Y => n98);
   U106 : NAND3X1 port map( A => n107, B => n108, C => n109, Y => n106);
   U107 : NAND3X1 port map( A => n110, B => n111, C => n112, Y => n108);
   U108 : NAND2X1 port map( A => n113, B => n114, Y => n111);
   U109 : AND2X2 port map( A => n117, B => n118, Y => n116);
   U110 : NAND2X1 port map( A => n21, B => n31, Y => n115);
   U111 : AND2X2 port map( A => n122, B => n123, Y => n113);
   U112 : XOR2X1 port map( A => B(16), B => A(16), Y => n104);
   U113 : NAND2X1 port map( A => n105, B => n109, Y => n125);
   U114 : OR2X2 port map( A => A(15), B => B(15), Y => n109);
   U115 : NAND2X1 port map( A => B(15), B => A(15), Y => n105);
   U116 : NAND2X1 port map( A => n112, B => n126, Y => n124);
   U117 : NAND2X1 port map( A => n127, B => n107, Y => n126);
   U118 : NAND2X1 port map( A => B(14), B => A(14), Y => n112);
   U119 : OR2X2 port map( A => A(14), B => B(14), Y => n107);
   U120 : OAI21X1 port map( A => n128, B => n129, C => n110, Y => n127);
   U121 : INVX2 port map( A => n130, Y => n129);
   U122 : INVX2 port map( A => n123, Y => n128);
   U123 : XNOR2X1 port map( A => n131, B => n130, Y => SUM(13));
   U124 : OAI21X1 port map( A => n132, B => n133, C => n117, Y => n130);
   U125 : INVX2 port map( A => n122, Y => n132);
   U126 : NAND2X1 port map( A => n123, B => n110, Y => n131);
   U127 : NAND2X1 port map( A => B(13), B => A(13), Y => n110);
   U128 : OR2X2 port map( A => A(13), B => B(13), Y => n123);
   U129 : NAND2X1 port map( A => B(12), B => A(12), Y => n117);
   U130 : OR2X2 port map( A => A(12), B => B(12), Y => n122);
   U131 : AND2X2 port map( A => n134, B => n118, Y => n133);
   U132 : NAND2X1 port map( A => n135, B => n136, Y => n118);
   U133 : NAND3X1 port map( A => n137, B => n138, C => n139, Y => n136);
   U134 : NAND3X1 port map( A => n29, B => n140, C => n141, Y => n138);
   U135 : NAND2X1 port map( A => n30, B => n33, Y => n140);
   U136 : NAND2X1 port map( A => n21, B => n31, Y => n134);
   U137 : NAND3X1 port map( A => n29, B => n34, C => n141, Y => n143);
   U138 : INVX2 port map( A => n135, Y => n142);
   U139 : NAND2X1 port map( A => n139, B => n135, Y => n145);
   U140 : OR2X2 port map( A => A(11), B => B(11), Y => n135);
   U141 : NAND2X1 port map( A => B(11), B => A(11), Y => n139);
   U142 : AOI21X1 port map( A => n146, B => n141, C => n147, Y => n144);
   U143 : NAND2X1 port map( A => B(10), B => A(10), Y => n137);
   U144 : OR2X2 port map( A => A(10), B => B(10), Y => n141);
   U145 : OAI21X1 port map( A => n28, B => n148, C => n30, Y => n146);
   U146 : NAND2X1 port map( A => B(9), B => A(9), Y => n30);
   U147 : INVX2 port map( A => n29, Y => n148);
   U148 : OR2X2 port map( A => A(9), B => B(9), Y => n29);
   U149 : AND2X2 port map( A => n149, B => n33, Y => n28);
   U150 : NAND2X1 port map( A => B(8), B => A(8), Y => n33);
   U151 : NAND2X1 port map( A => n34, B => n31, Y => n149);
   U152 : OAI21X1 port map( A => n119, B => n120, C => n121, Y => n31);
   U153 : NAND2X1 port map( A => n38, B => n150, Y => n121);
   U154 : NAND3X1 port map( A => n42, B => n151, C => n37, Y => n150);
   U155 : NAND2X1 port map( A => B(7), B => A(7), Y => n37);
   U156 : NAND3X1 port map( A => n46, B => n152, C => n40, Y => n151);
   U157 : NAND2X1 port map( A => n44, B => n48, Y => n152);
   U158 : NAND2X1 port map( A => B(4), B => A(4), Y => n48);
   U159 : NAND2X1 port map( A => B(5), B => A(5), Y => n44);
   U160 : NAND2X1 port map( A => B(6), B => A(6), Y => n42);
   U161 : OR2X2 port map( A => n153, B => n154, Y => n120);
   U162 : NAND3X1 port map( A => n46, B => n49, C => n40, Y => n154);
   U163 : OR2X2 port map( A => A(6), B => B(6), Y => n40);
   U164 : OR2X2 port map( A => A(4), B => B(4), Y => n49);
   U165 : OR2X2 port map( A => A(5), B => B(5), Y => n46);
   U166 : INVX2 port map( A => n38, Y => n153);
   U167 : OR2X2 port map( A => A(7), B => B(7), Y => n38);
   U168 : INVX2 port map( A => n155, Y => n119);
   U169 : OAI21X1 port map( A => n156, B => n157, C => n54, Y => n155);
   U170 : NAND2X1 port map( A => B(3), B => A(3), Y => n54);
   U171 : OAI21X1 port map( A => n158, B => n159, C => n53, Y => n157);
   U172 : OR2X2 port map( A => A(3), B => B(3), Y => n53);
   U173 : OAI21X1 port map( A => n160, B => n86, C => n58, Y => n159);
   U174 : NAND2X1 port map( A => B(2), B => A(2), Y => n58);
   U175 : INVX2 port map( A => n63, Y => n160);
   U176 : OR2X2 port map( A => A(1), B => B(1), Y => n63);
   U177 : INVX2 port map( A => n61, Y => n158);
   U178 : NAND2X1 port map( A => B(1), B => A(1), Y => n61);
   U179 : INVX2 port map( A => n56, Y => n156);
   U180 : OR2X2 port map( A => A(2), B => B(2), Y => n56);
   U181 : OR2X2 port map( A => A(8), B => B(8), Y => n34);
   U182 : NAND2X1 port map( A => B(0), B => A(0), Y => n86);
   U183 : OR2X2 port map( A => A(0), B => B(0), Y => n87);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW01_add_12 is

   port( A, B : in std_logic_vector (23 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (23 downto 0);  CO : out std_logic);

end matrix_math_DW01_add_12;

architecture SYN_cla of matrix_math_DW01_add_12 is

   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, SUM_19_port, 
      SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, SUM_14_port, 
      SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, n1, n2, 
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, SUM_8_port, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105 : std_logic;

begin
   SUM <= ( SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, SUM_19_port, 
      SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, SUM_14_port, 
      SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, B(7), B(6), B(5), B(4), B(3), B(2), B(1), B(0) );
   
   U2 : AND2X1 port map( A => n70, B => n63, Y => n69);
   U3 : AND2X2 port map( A => n94, B => n95, Y => n1);
   U4 : NAND2X1 port map( A => n30, B => A(16), Y => n2);
   U5 : OAI21X1 port map( A => n41, B => n42, C => n43, Y => n3);
   U6 : INVX1 port map( A => n53, Y => n4);
   U7 : INVX1 port map( A => n53, Y => n45);
   U8 : OR2X2 port map( A => n30, B => A(16), Y => n70);
   U9 : BUFX2 port map( A => B(16), Y => n30);
   U10 : OR2X2 port map( A => B(20), B => A(20), Y => n5);
   U11 : INVX1 port map( A => n5, Y => n6);
   U12 : INVX1 port map( A => n6, Y => n7);
   U13 : INVX1 port map( A => n13, Y => n8);
   U14 : INVX2 port map( A => n18, Y => n13);
   U15 : XOR2X1 port map( A => n54, B => n9, Y => SUM_20_port);
   U16 : NAND2X1 port map( A => n48, B => n5, Y => n9);
   U17 : NOR2X1 port map( A => B(22), B => A(22), Y => n10);
   U18 : INVX1 port map( A => n10, Y => n39);
   U19 : AND2X2 port map( A => B(22), B => A(22), Y => n26);
   U20 : BUFX4 port map( A => B(16), Y => n31);
   U21 : NAND2X1 port map( A => n2, B => n74, Y => n11);
   U22 : NAND2X1 port map( A => n11, B => n69, Y => n68);
   U23 : XOR2X1 port map( A => n50, B => n12, Y => SUM_21_port);
   U24 : AND2X2 port map( A => n44, B => n43, Y => n12);
   U25 : INVX1 port map( A => n8, Y => n62);
   U26 : INVX1 port map( A => B(18), Y => n14);
   U27 : INVX1 port map( A => n14, Y => n15);
   U28 : INVX1 port map( A => n17, Y => n16);
   U29 : AOI21X1 port map( A => n58, B => n57, C => n59, Y => n17);
   U30 : NOR2X1 port map( A => A(18), B => B(18), Y => n18);
   U31 : INVX1 port map( A => n96, Y => n104);
   U32 : AND2X1 port map( A => n31, B => A(16), Y => n28);
   U33 : AND2X1 port map( A => n32, B => n35, Y => SUM_8_port);
   U34 : XNOR2X1 port map( A => n67, B => n19, Y => SUM_18_port);
   U35 : NAND2X1 port map( A => n62, B => n61, Y => n19);
   U36 : XNOR2X1 port map( A => n45, B => n56, Y => SUM_19_port);
   U37 : XNOR2X1 port map( A => n89, B => n20, Y => SUM_14_port);
   U38 : NAND2X1 port map( A => n79, B => n90, Y => n20);
   U39 : XOR2X1 port map( A => n101, B => n102, Y => SUM_11_port);
   U40 : XOR2X1 port map( A => n91, B => n21, Y => SUM_13_port);
   U41 : NAND2X1 port map( A => n92, B => n82, Y => n21);
   U42 : XNOR2X1 port map( A => n1, B => n22, Y => SUM_12_port);
   U43 : NAND2X1 port map( A => n84, B => n85, Y => n22);
   U44 : XNOR2X1 port map( A => n103, B => n23, Y => SUM_10_port);
   U45 : NAND2X1 port map( A => n100, B => n96, Y => n23);
   U46 : XOR2X1 port map( A => n32, B => n24, Y => SUM_9_port);
   U47 : NAND2X1 port map( A => n33, B => n34, Y => n24);
   U48 : XOR2X1 port map( A => n71, B => n25, Y => SUM_17_port);
   U49 : NAND2X1 port map( A => n63, B => n60, Y => n25);
   U50 : NOR2X1 port map( A => A(15), B => B(15), Y => n27);
   U51 : OR2X1 port map( A => A(16), B => n31, Y => n72);
   U52 : XNOR2X1 port map( A => n36, B => n37, Y => SUM_23_port);
   U53 : XOR2X1 port map( A => B(23), B => A(23), Y => n37);
   U54 : AOI21X1 port map( A => n38, B => n39, C => n26, Y => n36);
   U55 : XOR2X1 port map( A => n40, B => n3, Y => SUM_22_port);
   U56 : NOR2X1 port map( A => n10, B => n26, Y => n40);
   U57 : OAI21X1 port map( A => n42, B => n41, C => n43, Y => n38);
   U58 : NAND2X1 port map( A => n7, B => n44, Y => n42);
   U59 : AOI21X1 port map( A => n4, B => n46, C => n47, Y => n41);
   U60 : NAND2X1 port map( A => n48, B => n49, Y => n47);
   U61 : OR2X2 port map( A => B(21), B => A(21), Y => n44);
   U62 : NAND2X1 port map( A => B(21), B => A(21), Y => n43);
   U63 : NAND2X1 port map( A => n48, B => n51, Y => n50);
   U64 : NAND3X1 port map( A => n46, B => n5, C => n52, Y => n51);
   U65 : NAND2X1 port map( A => n53, B => n49, Y => n52);
   U66 : NAND2X1 port map( A => B(20), B => A(20), Y => n48);
   U67 : AOI21X1 port map( A => n16, B => n46, C => n55, Y => n54);
   U68 : INVX2 port map( A => n49, Y => n55);
   U69 : NAND2X1 port map( A => n49, B => n46, Y => n56);
   U70 : OR2X2 port map( A => A(19), B => B(19), Y => n46);
   U71 : NAND2X1 port map( A => B(19), B => A(19), Y => n49);
   U72 : AOI21X1 port map( A => n58, B => n57, C => n59, Y => n53);
   U73 : OAI21X1 port map( A => n18, B => n60, C => n61, Y => n59);
   U74 : AND2X2 port map( A => n13, B => n63, Y => n58);
   U75 : AOI21X1 port map( A => n64, B => n74, C => n65, Y => n57);
   U76 : NOR2X1 port map( A => A(16), B => n31, Y => n65);
   U77 : NAND2X1 port map( A => n31, B => A(16), Y => n64);
   U78 : NAND2X1 port map( A => n15, B => A(18), Y => n61);
   U79 : NAND2X1 port map( A => n60, B => n68, Y => n67);
   U80 : NAND2X1 port map( A => B(17), B => A(17), Y => n60);
   U81 : OR2X2 port map( A => B(17), B => A(17), Y => n63);
   U82 : AOI21X1 port map( A => n66, B => n72, C => n28, Y => n71);
   U83 : XNOR2X1 port map( A => n73, B => n74, Y => SUM_16_port);
   U84 : INVX2 port map( A => n66, Y => n74);
   U85 : OAI21X1 port map( A => n27, B => n75, C => n76, Y => n66);
   U86 : OAI21X1 port map( A => n77, B => n78, C => n79, Y => n75);
   U87 : OAI21X1 port map( A => n80, B => n81, C => n82, Y => n78);
   U88 : OAI21X1 port map( A => n83, B => n1, C => n84, Y => n81);
   U89 : INVX2 port map( A => n85, Y => n83);
   U90 : XOR2X1 port map( A => n31, B => A(16), Y => n73);
   U91 : XNOR2X1 port map( A => n86, B => n87, Y => SUM_15_port);
   U92 : NOR2X1 port map( A => n88, B => n27, Y => n87);
   U93 : INVX2 port map( A => n76, Y => n88);
   U94 : NAND2X1 port map( A => B(15), B => A(15), Y => n76);
   U95 : AOI21X1 port map( A => n89, B => n79, C => n77, Y => n86);
   U96 : INVX2 port map( A => n90, Y => n77);
   U97 : NAND2X1 port map( A => B(14), B => A(14), Y => n90);
   U98 : OR2X2 port map( A => A(14), B => B(14), Y => n79);
   U99 : OAI21X1 port map( A => n80, B => n91, C => n82, Y => n89);
   U100 : INVX2 port map( A => n92, Y => n80);
   U101 : NAND2X1 port map( A => B(13), B => A(13), Y => n82);
   U102 : OR2X2 port map( A => A(13), B => B(13), Y => n92);
   U103 : AND2X2 port map( A => n93, B => n85, Y => n91);
   U104 : NAND2X1 port map( A => n1, B => n84, Y => n93);
   U105 : NAND2X1 port map( A => B(12), B => A(12), Y => n85);
   U106 : OR2X2 port map( A => A(12), B => B(12), Y => n84);
   U107 : NAND3X1 port map( A => n96, B => n97, C => n98, Y => n95);
   U108 : NAND3X1 port map( A => n33, B => n99, C => n100, Y => n97);
   U109 : NAND2X1 port map( A => n34, B => n32, Y => n99);
   U110 : NAND2X1 port map( A => n98, B => n94, Y => n102);
   U111 : OR2X2 port map( A => A(11), B => B(11), Y => n94);
   U112 : NAND2X1 port map( A => B(11), B => A(11), Y => n98);
   U113 : AOI21X1 port map( A => n103, B => n100, C => n104, Y => n101);
   U114 : NAND2X1 port map( A => B(10), B => A(10), Y => n96);
   U115 : OR2X2 port map( A => A(10), B => B(10), Y => n100);
   U116 : OAI21X1 port map( A => n32, B => n105, C => n34, Y => n103);
   U117 : NAND2X1 port map( A => B(9), B => A(9), Y => n34);
   U118 : INVX2 port map( A => n33, Y => n105);
   U119 : OR2X2 port map( A => A(9), B => B(9), Y => n33);
   U120 : NAND2X1 port map( A => B(8), B => A(8), Y => n32);
   U121 : OR2X2 port map( A => A(8), B => B(8), Y => n35);

end SYN_cla;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW02_mult_2 is

   port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  PRODUCT
         : out std_logic_vector (31 downto 0));

end matrix_math_DW02_mult_2;

architecture SYN_csa of matrix_math_DW02_mult_2 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component matrix_math_DW01_add_25
      port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (29 downto 0);  CO : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_15_15_port, ab_15_14_port, ab_15_13_port, 
      ab_15_12_port, ab_15_11_port, ab_15_10_port, ab_15_9_port, ab_15_8_port, 
      ab_15_7_port, ab_15_6_port, ab_15_5_port, ab_15_4_port, ab_15_3_port, 
      ab_15_2_port, ab_15_1_port, ab_15_0_port, ab_14_15_port, ab_14_14_port, 
      ab_14_13_port, ab_14_12_port, ab_14_11_port, ab_14_10_port, ab_14_9_port,
      ab_14_8_port, ab_14_7_port, ab_14_6_port, ab_14_5_port, ab_14_4_port, 
      ab_14_3_port, ab_14_2_port, ab_14_1_port, ab_14_0_port, ab_13_15_port, 
      ab_13_14_port, ab_13_13_port, ab_13_12_port, ab_13_11_port, ab_13_10_port
      , ab_13_9_port, ab_13_8_port, ab_13_7_port, ab_13_6_port, ab_13_5_port, 
      ab_13_4_port, ab_13_3_port, ab_13_2_port, ab_13_1_port, ab_13_0_port, 
      ab_12_15_port, ab_12_14_port, ab_12_13_port, ab_12_12_port, ab_12_11_port
      , ab_12_10_port, ab_12_9_port, ab_12_8_port, ab_12_7_port, ab_12_6_port, 
      ab_12_5_port, ab_12_4_port, ab_12_3_port, ab_12_2_port, ab_12_1_port, 
      ab_12_0_port, ab_11_15_port, ab_11_14_port, ab_11_13_port, ab_11_12_port,
      ab_11_11_port, ab_11_10_port, ab_11_9_port, ab_11_8_port, ab_11_7_port, 
      ab_11_6_port, ab_11_5_port, ab_11_4_port, ab_11_3_port, ab_11_2_port, 
      ab_11_1_port, ab_11_0_port, ab_10_15_port, ab_10_14_port, ab_10_13_port, 
      ab_10_12_port, ab_10_11_port, ab_10_10_port, ab_10_9_port, ab_10_8_port, 
      ab_10_7_port, ab_10_6_port, ab_10_5_port, ab_10_4_port, ab_10_3_port, 
      ab_10_2_port, ab_10_1_port, ab_10_0_port, ab_9_15_port, ab_9_14_port, 
      ab_9_13_port, ab_9_12_port, ab_9_11_port, ab_9_10_port, ab_9_9_port, 
      ab_9_8_port, ab_9_7_port, ab_9_6_port, ab_9_5_port, ab_9_4_port, 
      ab_9_3_port, ab_9_2_port, ab_9_1_port, ab_9_0_port, ab_8_15_port, 
      ab_8_14_port, ab_8_13_port, ab_8_12_port, ab_8_11_port, ab_8_10_port, 
      ab_8_9_port, ab_8_8_port, ab_8_7_port, ab_8_6_port, ab_8_5_port, 
      ab_8_4_port, ab_8_3_port, ab_8_2_port, ab_8_1_port, ab_8_0_port, 
      ab_7_15_port, ab_7_14_port, ab_7_13_port, ab_7_12_port, ab_7_11_port, 
      ab_7_10_port, ab_7_9_port, ab_7_8_port, ab_7_7_port, ab_7_6_port, 
      ab_7_5_port, ab_7_4_port, ab_7_3_port, ab_7_2_port, ab_7_1_port, 
      ab_7_0_port, ab_6_15_port, ab_6_14_port, ab_6_13_port, ab_6_12_port, 
      ab_6_11_port, ab_6_10_port, ab_6_9_port, ab_6_8_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_15_port, ab_5_14_port, ab_5_13_port, 
      ab_5_12_port, ab_5_11_port, ab_5_10_port, ab_5_9_port, ab_5_8_port, 
      ab_5_7_port, ab_5_6_port, ab_5_5_port, ab_5_4_port, ab_5_3_port, 
      ab_5_2_port, ab_5_1_port, ab_5_0_port, ab_4_15_port, ab_4_14_port, 
      ab_4_13_port, ab_4_12_port, ab_4_11_port, ab_4_10_port, ab_4_9_port, 
      ab_4_8_port, ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, 
      ab_4_3_port, ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_15_port, 
      ab_3_14_port, ab_3_13_port, ab_3_12_port, ab_3_11_port, ab_3_10_port, 
      ab_3_9_port, ab_3_7_port, ab_3_6_port, ab_3_5_port, ab_3_4_port, 
      ab_3_3_port, ab_3_2_port, ab_3_1_port, ab_3_0_port, ab_2_15_port, 
      ab_2_14_port, ab_2_13_port, ab_2_12_port, ab_2_11_port, ab_2_10_port, 
      ab_2_9_port, ab_2_8_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, 
      ab_2_4_port, ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, 
      ab_1_15_port, ab_1_14_port, ab_1_12_port, ab_1_11_port, ab_1_10_port, 
      ab_1_9_port, ab_1_8_port, ab_1_7_port, ab_1_6_port, ab_1_5_port, 
      ab_1_4_port, ab_1_3_port, ab_1_2_port, ab_1_1_port, ab_1_0_port, 
      ab_0_14_port, ab_0_13_port, ab_0_12_port, ab_0_10_port, ab_0_9_port, 
      ab_0_8_port, ab_0_7_port, ab_0_6_port, ab_0_4_port, ab_0_3_port, 
      ab_0_2_port, ab_0_1_port, CARRYB_15_15_port, CARRYB_15_14_port, 
      CARRYB_15_13_port, CARRYB_15_12_port, CARRYB_15_11_port, 
      CARRYB_15_10_port, CARRYB_15_9_port, CARRYB_15_8_port, CARRYB_15_7_port, 
      CARRYB_15_6_port, CARRYB_15_5_port, CARRYB_15_4_port, CARRYB_15_3_port, 
      CARRYB_15_2_port, CARRYB_15_1_port, CARRYB_15_0_port, CARRYB_14_14_port, 
      CARRYB_14_13_port, CARRYB_14_12_port, CARRYB_14_11_port, 
      CARRYB_14_10_port, CARRYB_14_9_port, CARRYB_14_8_port, CARRYB_14_7_port, 
      CARRYB_14_6_port, CARRYB_14_5_port, CARRYB_14_4_port, CARRYB_14_3_port, 
      CARRYB_14_2_port, CARRYB_14_1_port, CARRYB_14_0_port, CARRYB_13_14_port, 
      CARRYB_13_13_port, CARRYB_13_12_port, CARRYB_13_11_port, 
      CARRYB_13_10_port, CARRYB_13_9_port, CARRYB_13_8_port, CARRYB_13_7_port, 
      CARRYB_13_6_port, CARRYB_13_4_port, CARRYB_13_2_port, CARRYB_13_1_port, 
      CARRYB_13_0_port, CARRYB_12_14_port, CARRYB_12_13_port, CARRYB_12_12_port
      , CARRYB_12_11_port, CARRYB_12_10_port, CARRYB_12_9_port, 
      CARRYB_12_8_port, CARRYB_12_7_port, CARRYB_12_6_port, CARRYB_12_5_port, 
      CARRYB_12_4_port, CARRYB_12_3_port, CARRYB_12_2_port, CARRYB_12_1_port, 
      CARRYB_12_0_port, CARRYB_11_14_port, CARRYB_11_13_port, CARRYB_11_12_port
      , CARRYB_11_11_port, CARRYB_11_10_port, CARRYB_11_9_port, 
      CARRYB_11_8_port, CARRYB_11_7_port, CARRYB_11_6_port, CARRYB_11_5_port, 
      CARRYB_11_4_port, CARRYB_11_3_port, CARRYB_11_2_port, CARRYB_11_1_port, 
      CARRYB_11_0_port, CARRYB_10_14_port, CARRYB_10_13_port, CARRYB_10_12_port
      , CARRYB_10_11_port, CARRYB_10_10_port, CARRYB_10_9_port, 
      CARRYB_10_8_port, CARRYB_10_7_port, CARRYB_10_6_port, CARRYB_10_5_port, 
      CARRYB_10_4_port, CARRYB_10_3_port, CARRYB_10_2_port, CARRYB_10_1_port, 
      CARRYB_10_0_port, CARRYB_9_14_port, CARRYB_9_13_port, CARRYB_9_12_port, 
      CARRYB_9_11_port, CARRYB_9_10_port, CARRYB_9_9_port, CARRYB_9_8_port, 
      CARRYB_9_7_port, CARRYB_9_6_port, CARRYB_9_5_port, CARRYB_9_4_port, 
      CARRYB_9_3_port, CARRYB_9_2_port, CARRYB_9_1_port, CARRYB_9_0_port, 
      CARRYB_8_14_port, CARRYB_8_13_port, CARRYB_8_12_port, CARRYB_8_11_port, 
      CARRYB_8_10_port, CARRYB_8_9_port, CARRYB_8_8_port, CARRYB_8_7_port, 
      CARRYB_8_6_port, CARRYB_8_5_port, CARRYB_8_4_port, CARRYB_8_3_port, 
      CARRYB_8_2_port, CARRYB_8_1_port, CARRYB_8_0_port, CARRYB_7_14_port, 
      CARRYB_7_13_port, CARRYB_7_12_port, CARRYB_7_11_port, CARRYB_7_10_port, 
      CARRYB_7_9_port, CARRYB_7_8_port, CARRYB_7_7_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_14_port, CARRYB_6_13_port, 
      CARRYB_6_12_port, CARRYB_6_11_port, CARRYB_6_10_port, CARRYB_6_9_port, 
      CARRYB_6_8_port, CARRYB_6_7_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_14_port, CARRYB_5_13_port, CARRYB_5_12_port, 
      CARRYB_5_10_port, CARRYB_5_9_port, CARRYB_5_8_port, CARRYB_5_7_port, 
      CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, CARRYB_5_3_port, 
      CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, CARRYB_4_14_port, 
      CARRYB_4_13_port, CARRYB_4_12_port, CARRYB_4_11_port, CARRYB_4_9_port, 
      CARRYB_4_8_port, CARRYB_4_7_port, CARRYB_4_6_port, CARRYB_4_5_port, 
      CARRYB_4_4_port, CARRYB_4_3_port, CARRYB_4_2_port, CARRYB_4_1_port, 
      CARRYB_4_0_port, CARRYB_3_14_port, CARRYB_3_13_port, CARRYB_3_12_port, 
      CARRYB_3_11_port, CARRYB_3_10_port, CARRYB_3_9_port, CARRYB_3_8_port, 
      CARRYB_3_7_port, CARRYB_3_6_port, CARRYB_3_5_port, CARRYB_3_4_port, 
      CARRYB_3_3_port, CARRYB_3_2_port, CARRYB_3_1_port, CARRYB_3_0_port, 
      CARRYB_2_14_port, CARRYB_2_13_port, CARRYB_2_12_port, CARRYB_2_11_port, 
      CARRYB_2_10_port, CARRYB_2_9_port, CARRYB_2_7_port, CARRYB_2_6_port, 
      CARRYB_2_5_port, CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, 
      CARRYB_2_1_port, CARRYB_2_0_port, CARRYB_1_1_port, SUMB_15_15_port, 
      SUMB_15_14_port, SUMB_15_13_port, SUMB_15_12_port, SUMB_15_11_port, 
      SUMB_15_10_port, SUMB_15_9_port, SUMB_15_8_port, SUMB_15_7_port, 
      SUMB_15_6_port, SUMB_15_5_port, SUMB_15_4_port, SUMB_15_3_port, 
      SUMB_15_2_port, SUMB_15_1_port, SUMB_15_0_port, SUMB_14_14_port, 
      SUMB_14_13_port, SUMB_14_12_port, SUMB_14_11_port, SUMB_14_10_port, 
      SUMB_14_9_port, SUMB_14_8_port, SUMB_14_7_port, SUMB_14_6_port, 
      SUMB_14_5_port, SUMB_14_4_port, SUMB_14_3_port, SUMB_14_2_port, 
      SUMB_14_1_port, SUMB_13_14_port, SUMB_13_13_port, SUMB_13_12_port, 
      SUMB_13_11_port, SUMB_13_10_port, SUMB_13_9_port, SUMB_13_8_port, 
      SUMB_13_7_port, SUMB_13_6_port, SUMB_13_5_port, SUMB_13_4_port, 
      SUMB_13_3_port, SUMB_13_2_port, SUMB_13_1_port, SUMB_12_14_port, 
      SUMB_12_13_port, SUMB_12_12_port, SUMB_12_11_port, SUMB_12_10_port, 
      SUMB_12_9_port, SUMB_12_8_port, SUMB_12_7_port, SUMB_12_6_port, 
      SUMB_12_5_port, SUMB_12_4_port, SUMB_12_3_port, SUMB_12_2_port, 
      SUMB_12_1_port, SUMB_11_14_port, SUMB_11_13_port, SUMB_11_12_port, 
      SUMB_11_11_port, SUMB_11_10_port, SUMB_11_9_port, SUMB_11_8_port, 
      SUMB_11_7_port, SUMB_11_6_port, SUMB_11_5_port, SUMB_11_4_port, 
      SUMB_11_3_port, SUMB_11_2_port, SUMB_11_1_port, SUMB_10_14_port, 
      SUMB_10_13_port, SUMB_10_12_port, SUMB_10_11_port, SUMB_10_10_port, 
      SUMB_10_9_port, SUMB_10_8_port, SUMB_10_7_port, SUMB_10_6_port, 
      SUMB_10_5_port, SUMB_10_4_port, SUMB_10_3_port, SUMB_10_2_port, 
      SUMB_10_1_port, SUMB_9_14_port, SUMB_9_13_port, SUMB_9_12_port, 
      SUMB_9_11_port, SUMB_9_10_port, SUMB_9_9_port, SUMB_9_8_port, 
      SUMB_9_7_port, SUMB_9_6_port, SUMB_9_5_port, SUMB_9_4_port, SUMB_9_3_port
      , SUMB_9_2_port, SUMB_9_1_port, SUMB_8_14_port, SUMB_8_13_port, 
      SUMB_8_12_port, SUMB_8_11_port, SUMB_8_10_port, SUMB_8_9_port, 
      SUMB_8_8_port, SUMB_8_7_port, SUMB_8_6_port, SUMB_8_5_port, SUMB_8_4_port
      , SUMB_8_3_port, SUMB_8_2_port, SUMB_8_1_port, SUMB_7_14_port, 
      SUMB_7_13_port, SUMB_7_12_port, SUMB_7_11_port, SUMB_7_10_port, 
      SUMB_7_9_port, SUMB_7_8_port, SUMB_7_7_port, SUMB_7_6_port, SUMB_7_5_port
      , SUMB_7_4_port, SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, 
      SUMB_6_14_port, SUMB_6_13_port, SUMB_6_12_port, SUMB_6_11_port, 
      SUMB_6_10_port, SUMB_6_9_port, SUMB_6_8_port, SUMB_6_7_port, 
      SUMB_6_6_port, SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port
      , SUMB_6_1_port, SUMB_5_14_port, SUMB_5_13_port, SUMB_5_12_port, 
      SUMB_5_11_port, SUMB_5_10_port, SUMB_5_9_port, SUMB_5_8_port, 
      SUMB_5_7_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_14_port, SUMB_4_13_port, 
      SUMB_4_12_port, SUMB_4_11_port, SUMB_4_10_port, SUMB_4_9_port, 
      SUMB_4_8_port, SUMB_4_7_port, SUMB_4_6_port, SUMB_4_5_port, SUMB_4_4_port
      , SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_14_port, 
      SUMB_3_13_port, SUMB_3_12_port, SUMB_3_11_port, SUMB_3_10_port, 
      SUMB_3_9_port, SUMB_3_8_port, SUMB_3_7_port, SUMB_3_6_port, SUMB_3_5_port
      , SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, SUMB_3_1_port, 
      SUMB_2_14_port, SUMB_2_13_port, SUMB_2_12_port, SUMB_2_11_port, 
      SUMB_2_10_port, SUMB_2_9_port, SUMB_2_8_port, SUMB_2_7_port, 
      SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port, SUMB_2_2_port
      , SUMB_2_1_port, SUMB_1_14_port, SUMB_1_13_port, SUMB_1_12_port, 
      SUMB_1_11_port, SUMB_1_10_port, SUMB_1_9_port, SUMB_1_8_port, 
      SUMB_1_7_port, SUMB_1_6_port, SUMB_1_5_port, SUMB_1_4_port, SUMB_1_3_port
      , SUMB_1_2_port, SUMB_1_1_port, A1_28_port, A1_27_port, A1_26_port, 
      A1_25_port, A1_24_port, A1_23_port, A1_22_port, A1_21_port, A1_20_port, 
      A1_19_port, A1_18_port, A1_17_port, A1_16_port, A1_15_port, A1_14_port, 
      A1_13_port, A1_12_port, A1_11_port, A1_10_port, A1_9_port, A1_8_port, 
      A1_7_port, A1_6_port, A1_5_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, A2_22_port, A2_21_port, A2_14_port, n3, n4, n5, n6,
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, 
      n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, 
      n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_8 : FAX1 port map( A => ab_15_8_port, B => CARRYB_14_8_port, C => 
                           SUMB_14_9_port, YC => CARRYB_15_8_port, YS => 
                           SUMB_15_8_port);
   S4_9 : FAX1 port map( A => ab_15_9_port, B => CARRYB_14_9_port, C => 
                           SUMB_14_10_port, YC => CARRYB_15_9_port, YS => 
                           SUMB_15_9_port);
   S4_10 : FAX1 port map( A => ab_15_10_port, B => CARRYB_14_10_port, C => 
                           SUMB_14_11_port, YC => CARRYB_15_10_port, YS => 
                           SUMB_15_10_port);
   S4_11 : FAX1 port map( A => ab_15_11_port, B => CARRYB_14_11_port, C => 
                           SUMB_14_12_port, YC => CARRYB_15_11_port, YS => 
                           SUMB_15_11_port);
   S4_12 : FAX1 port map( A => ab_15_12_port, B => CARRYB_14_12_port, C => 
                           SUMB_14_13_port, YC => CARRYB_15_12_port, YS => 
                           SUMB_15_12_port);
   S4_13 : FAX1 port map( A => ab_15_13_port, B => CARRYB_14_13_port, C => 
                           SUMB_14_14_port, YC => CARRYB_15_13_port, YS => 
                           SUMB_15_13_port);
   S5_14 : FAX1 port map( A => ab_15_14_port, B => CARRYB_14_14_port, C => 
                           ab_14_15_port, YC => CARRYB_15_14_port, YS => 
                           SUMB_15_14_port);
   S14_15 : FAX1 port map( A => n1052, B => n1051, C => ab_15_15_port, YC => 
                           CARRYB_15_15_port, YS => SUMB_15_15_port);
   S2_14_9 : FAX1 port map( A => ab_14_9_port, B => CARRYB_13_9_port, C => 
                           SUMB_13_10_port, YC => CARRYB_14_9_port, YS => 
                           SUMB_14_9_port);
   S2_14_10 : FAX1 port map( A => ab_14_10_port, B => CARRYB_13_10_port, C => 
                           SUMB_13_11_port, YC => CARRYB_14_10_port, YS => 
                           SUMB_14_10_port);
   S2_14_11 : FAX1 port map( A => ab_14_11_port, B => CARRYB_13_11_port, C => 
                           SUMB_13_12_port, YC => CARRYB_14_11_port, YS => 
                           SUMB_14_11_port);
   S2_14_12 : FAX1 port map( A => ab_14_12_port, B => CARRYB_13_12_port, C => 
                           SUMB_13_13_port, YC => CARRYB_14_12_port, YS => 
                           SUMB_14_12_port);
   S2_14_13 : FAX1 port map( A => ab_14_13_port, B => CARRYB_13_13_port, C => 
                           SUMB_13_14_port, YC => CARRYB_14_13_port, YS => 
                           SUMB_14_13_port);
   S3_14_14 : FAX1 port map( A => ab_14_14_port, B => CARRYB_13_14_port, C => 
                           ab_13_15_port, YC => CARRYB_14_14_port, YS => 
                           SUMB_14_14_port);
   S2_13_9 : FAX1 port map( A => ab_13_9_port, B => CARRYB_12_9_port, C => 
                           SUMB_12_10_port, YC => CARRYB_13_9_port, YS => 
                           SUMB_13_9_port);
   S2_13_10 : FAX1 port map( A => ab_13_10_port, B => CARRYB_12_10_port, C => 
                           SUMB_12_11_port, YC => CARRYB_13_10_port, YS => 
                           SUMB_13_10_port);
   S2_13_11 : FAX1 port map( A => ab_13_11_port, B => CARRYB_12_11_port, C => 
                           SUMB_12_12_port, YC => CARRYB_13_11_port, YS => 
                           SUMB_13_11_port);
   S2_13_12 : FAX1 port map( A => ab_13_12_port, B => CARRYB_12_12_port, C => 
                           SUMB_12_13_port, YC => CARRYB_13_12_port, YS => 
                           SUMB_13_12_port);
   S2_13_13 : FAX1 port map( A => ab_13_13_port, B => CARRYB_12_13_port, C => 
                           SUMB_12_14_port, YC => CARRYB_13_13_port, YS => 
                           SUMB_13_13_port);
   S3_13_14 : FAX1 port map( A => ab_13_14_port, B => CARRYB_12_14_port, C => 
                           ab_12_15_port, YC => CARRYB_13_14_port, YS => 
                           SUMB_13_14_port);
   S2_12_11 : FAX1 port map( A => ab_12_11_port, B => CARRYB_11_11_port, C => 
                           SUMB_11_12_port, YC => CARRYB_12_11_port, YS => 
                           SUMB_12_11_port);
   S2_12_12 : FAX1 port map( A => ab_12_12_port, B => CARRYB_11_12_port, C => 
                           SUMB_11_13_port, YC => CARRYB_12_12_port, YS => 
                           SUMB_12_12_port);
   S2_12_13 : FAX1 port map( A => ab_12_13_port, B => CARRYB_11_13_port, C => 
                           SUMB_11_14_port, YC => CARRYB_12_13_port, YS => 
                           SUMB_12_13_port);
   S3_12_14 : FAX1 port map( A => ab_12_14_port, B => CARRYB_11_14_port, C => 
                           ab_11_15_port, YC => CARRYB_12_14_port, YS => 
                           SUMB_12_14_port);
   S2_11_1 : FAX1 port map( A => ab_11_1_port, B => CARRYB_10_1_port, C => 
                           SUMB_10_2_port, YC => CARRYB_11_1_port, YS => 
                           SUMB_11_1_port);
   S2_11_9 : FAX1 port map( A => ab_11_9_port, B => CARRYB_10_9_port, C => 
                           SUMB_10_10_port, YC => CARRYB_11_9_port, YS => 
                           SUMB_11_9_port);
   S2_11_12 : FAX1 port map( A => ab_11_12_port, B => CARRYB_10_12_port, C => 
                           SUMB_10_13_port, YC => CARRYB_11_12_port, YS => 
                           SUMB_11_12_port);
   S2_11_13 : FAX1 port map( A => ab_11_13_port, B => CARRYB_10_13_port, C => 
                           SUMB_10_14_port, YC => CARRYB_11_13_port, YS => 
                           SUMB_11_13_port);
   S3_11_14 : FAX1 port map( A => ab_11_14_port, B => CARRYB_10_14_port, C => 
                           ab_10_15_port, YC => CARRYB_11_14_port, YS => 
                           SUMB_11_14_port);
   S2_10_12 : FAX1 port map( A => ab_10_12_port, B => CARRYB_9_12_port, C => 
                           SUMB_9_13_port, YC => CARRYB_10_12_port, YS => 
                           SUMB_10_12_port);
   S2_10_13 : FAX1 port map( A => ab_10_13_port, B => CARRYB_9_13_port, C => 
                           SUMB_9_14_port, YC => CARRYB_10_13_port, YS => 
                           SUMB_10_13_port);
   S3_10_14 : FAX1 port map( A => ab_10_14_port, B => CARRYB_9_14_port, C => 
                           ab_9_15_port, YC => CARRYB_10_14_port, YS => 
                           SUMB_10_14_port);
   S1_9_0 : FAX1 port map( A => ab_9_0_port, B => CARRYB_8_0_port, C => 
                           SUMB_8_1_port, YC => CARRYB_9_0_port, YS => 
                           A1_7_port);
   S2_9_13 : FAX1 port map( A => ab_9_13_port, B => CARRYB_8_13_port, C => 
                           SUMB_8_14_port, YC => CARRYB_9_13_port, YS => 
                           SUMB_9_13_port);
   S3_9_14 : FAX1 port map( A => ab_9_14_port, B => CARRYB_8_14_port, C => 
                           ab_8_15_port, YC => CARRYB_9_14_port, YS => 
                           SUMB_9_14_port);
   S2_8_13 : FAX1 port map( A => ab_8_13_port, B => SUMB_7_14_port, C => 
                           CARRYB_7_13_port, YC => CARRYB_8_13_port, YS => 
                           SUMB_8_13_port);
   S3_8_14 : FAX1 port map( A => ab_8_14_port, B => CARRYB_7_14_port, C => 
                           ab_7_15_port, YC => CARRYB_8_14_port, YS => 
                           SUMB_8_14_port);
   S3_7_14 : FAX1 port map( A => ab_7_14_port, B => CARRYB_6_14_port, C => 
                           ab_6_15_port, YC => CARRYB_7_14_port, YS => 
                           SUMB_7_14_port);
   S1_6_0 : FAX1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, C => 
                           SUMB_5_1_port, YC => CARRYB_6_0_port, YS => 
                           A1_4_port);
   S2_6_1 : FAX1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, C => 
                           SUMB_5_2_port, YC => CARRYB_6_1_port, YS => 
                           SUMB_6_1_port);
   S2_6_12 : FAX1 port map( A => ab_6_12_port, B => n286, C => SUMB_5_13_port, 
                           YC => CARRYB_6_12_port, YS => SUMB_6_12_port);
   S2_6_13 : FAX1 port map( A => ab_6_13_port, B => n242, C => SUMB_5_14_port, 
                           YC => CARRYB_6_13_port, YS => SUMB_6_13_port);
   S2_5_12 : FAX1 port map( A => ab_5_12_port, B => CARRYB_4_12_port, C => 
                           SUMB_4_13_port, YC => CARRYB_5_12_port, YS => 
                           SUMB_5_12_port);
   S2_5_13 : FAX1 port map( A => ab_5_13_port, B => n367, C => SUMB_4_14_port, 
                           YC => CARRYB_5_13_port, YS => SUMB_5_13_port);
   S3_5_14 : FAX1 port map( A => ab_5_14_port, B => CARRYB_4_14_port, C => 
                           ab_4_15_port, YC => CARRYB_5_14_port, YS => 
                           SUMB_5_14_port);
   S1_4_0 : FAX1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, C => 
                           SUMB_3_1_port, YC => CARRYB_4_0_port, YS => 
                           A1_2_port);
   S2_4_13 : FAX1 port map( A => ab_4_13_port, B => CARRYB_3_13_port, C => 
                           SUMB_3_14_port, YC => CARRYB_4_13_port, YS => 
                           SUMB_4_13_port);
   S1_3_0 : FAX1 port map( A => ab_3_0_port, B => n968, C => SUMB_2_1_port, YC 
                           => CARRYB_3_0_port, YS => A1_1_port);
   S1_2_0 : FAX1 port map( A => ab_2_0_port, B => n958, C => SUMB_1_1_port, YC 
                           => CARRYB_2_0_port, YS => A1_0_port);
   S2_2_1 : FAX1 port map( A => ab_2_1_port, B => CARRYB_1_1_port, C => 
                           SUMB_1_2_port, YC => CARRYB_2_1_port, YS => 
                           SUMB_2_1_port);
   FS_1 : matrix_math_DW01_add_25 port map( A(29) => n1050, A(28) => A1_28_port
                           , A(27) => A1_27_port, A(26) => A1_26_port, A(25) =>
                           A1_25_port, A(24) => A1_24_port, A(23) => A1_23_port
                           , A(22) => A1_22_port, A(21) => A1_21_port, A(20) =>
                           A1_20_port, A(19) => A1_19_port, A(18) => A1_18_port
                           , A(17) => A1_17_port, A(16) => A1_16_port, A(15) =>
                           A1_15_port, A(14) => A1_14_port, A(13) => A1_13_port
                           , A(12) => A1_12_port, A(11) => A1_11_port, A(10) =>
                           A1_10_port, A(9) => A1_9_port, A(8) => A1_8_port, 
                           A(7) => A1_7_port, A(6) => A1_6_port, A(5) => 
                           A1_5_port, A(4) => A1_4_port, A(3) => A1_3_port, 
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(29) => n72, B(28) => n71, B(27) => n70,
                           B(26) => n69, B(25) => n68, B(24) => n67, B(23) => 
                           n66, B(22) => A2_22_port, B(21) => A2_21_port, B(20)
                           => n957, B(19) => n956, B(18) => n954, B(17) => n952
                           , B(16) => n953, B(15) => n955, B(14) => A2_14_port,
                           B(13) => n1055, B(12) => n1055, B(11) => n1055, 
                           B(10) => n1055, B(9) => n1055, B(8) => n1055, B(7) 
                           => n1055, B(6) => n1055, B(5) => n1055, B(4) => 
                           n1055, B(3) => n1055, B(2) => n1055, B(1) => n1055, 
                           B(0) => X_Logic0_port, CI => X_Logic0_port, SUM(29) 
                           => n_1159, SUM(28) => n_1160, SUM(27) => n_1161, 
                           SUM(26) => n_1162, SUM(25) => n_1163, SUM(24) => 
                           n_1164, SUM(23) => n_1165, SUM(22) => n_1166, 
                           SUM(21) => PRODUCT(23), SUM(20) => PRODUCT(22), 
                           SUM(19) => PRODUCT(21), SUM(18) => PRODUCT(20), 
                           SUM(17) => PRODUCT(19), SUM(16) => PRODUCT(18), 
                           SUM(15) => PRODUCT(17), SUM(14) => PRODUCT(16), 
                           SUM(13) => PRODUCT(15), SUM(12) => PRODUCT(14), 
                           SUM(11) => PRODUCT(13), SUM(10) => PRODUCT(12), 
                           SUM(9) => PRODUCT(11), SUM(8) => PRODUCT(10), SUM(7)
                           => PRODUCT(9), SUM(6) => PRODUCT(8), SUM(5) => 
                           PRODUCT(7), SUM(4) => PRODUCT(6), SUM(3) => 
                           PRODUCT(5), SUM(2) => PRODUCT(4), SUM(1) => 
                           PRODUCT(3), SUM(0) => PRODUCT(2), CO => n_1167);
   U2 : XOR2X1 port map( A => n3, B => ab_0_10_port, Y => SUMB_1_9_port);
   U3 : AND2X2 port map( A => n423, B => B(9), Y => n3);
   U4 : INVX2 port map( A => n1019, Y => n4);
   U5 : INVX2 port map( A => n1019, Y => n5);
   U6 : INVX2 port map( A => n1019, Y => n1020);
   U7 : INVX2 port map( A => A(2), Y => n1019);
   U8 : INVX4 port map( A => n1017, Y => n423);
   U9 : INVX1 port map( A => SUMB_2_7_port, Y => n323);
   U10 : XNOR2X1 port map( A => n282, B => n41, Y => n6);
   U11 : INVX2 port map( A => n8, Y => n9);
   U12 : NAND3X1 port map( A => n259, B => n258, C => n260, Y => n7);
   U13 : INVX1 port map( A => n1018, Y => n8);
   U14 : BUFX2 port map( A => n5, Y => n10);
   U15 : NAND3X1 port map( A => n335, B => n336, C => n337, Y => n11);
   U16 : BUFX2 port map( A => n418, Y => n12);
   U17 : XOR2X1 port map( A => CARRYB_6_6_port, B => n13, Y => n19);
   U18 : INVX8 port map( A => ab_7_6_port, Y => n13);
   U19 : NAND3X1 port map( A => n511, B => n510, C => n509, Y => n14);
   U20 : NAND3X1 port map( A => n455, B => n454, C => n456, Y => n15);
   U21 : XOR2X1 port map( A => n16, B => n373, Y => SUMB_8_4_port);
   U22 : INVX1 port map( A => SUMB_7_5_port, Y => n16);
   U23 : XNOR2X1 port map( A => n17, B => SUMB_4_7_port, Y => SUMB_5_6_port);
   U24 : XNOR2X1 port map( A => CARRYB_4_6_port, B => ab_5_6_port, Y => n17);
   U25 : BUFX2 port map( A => SUMB_5_11_port, Y => n18);
   U26 : INVX2 port map( A => A(0), Y => n1016);
   U27 : XOR2X1 port map( A => n374, B => n19, Y => SUMB_7_6_port);
   U28 : NAND3X1 port map( A => n746, B => n747, C => n748, Y => n20);
   U29 : AND2X1 port map( A => n423, B => B(9), Y => ab_1_9_port);
   U30 : INVX1 port map( A => SUMB_14_6_port, Y => n21);
   U31 : INVX1 port map( A => n21, Y => n22);
   U32 : XOR2X1 port map( A => CARRYB_13_2_port, B => n23, Y => n315);
   U33 : INVX8 port map( A => ab_14_2_port, Y => n23);
   U34 : XNOR2X1 port map( A => n24, B => n174, Y => SUMB_4_5_port);
   U35 : XOR2X1 port map( A => n407, B => ab_4_5_port, Y => n24);
   U36 : XNOR2X1 port map( A => CARRYB_14_0_port, B => n25, Y => n302);
   U37 : INVX8 port map( A => ab_15_0_port, Y => n25);
   U38 : BUFX4 port map( A => ab_2_12_port, Y => n160);
   U39 : XOR2X1 port map( A => SUMB_15_3_port, B => CARRYB_15_2_port, Y => 
                           A1_16_port);
   U40 : INVX1 port map( A => CARRYB_15_2_port, Y => n593);
   U41 : XNOR2X1 port map( A => n26, B => n347, Y => SUMB_10_2_port);
   U42 : XOR2X1 port map( A => CARRYB_9_2_port, B => ab_10_2_port, Y => n26);
   U43 : XOR2X1 port map( A => n134, B => n27, Y => n504);
   U44 : INVX8 port map( A => ab_14_3_port, Y => n27);
   U45 : XOR2X1 port map( A => n229, B => n29, Y => n28);
   U46 : XOR2X1 port map( A => n229, B => n29, Y => SUMB_12_3_port);
   U47 : AND2X2 port map( A => n766, B => n102, Y => n29);
   U48 : AND2X2 port map( A => n984, B => ab_1_14_port, Y => n30);
   U49 : XNOR2X1 port map( A => n31, B => CARRYB_11_8_port, Y => n642);
   U50 : INVX8 port map( A => ab_12_8_port, Y => n31);
   U51 : AND2X1 port map( A => SUMB_15_6_port, B => CARRYB_15_5_port, Y => n957
                           );
   U52 : XNOR2X1 port map( A => n32, B => n33, Y => SUMB_9_5_port);
   U53 : XNOR2X1 port map( A => CARRYB_8_5_port, B => ab_9_5_port, Y => n32);
   U54 : XOR2X1 port map( A => n447, B => n448, Y => n33);
   U55 : XOR2X1 port map( A => n34, B => SUMB_10_7_port, Y => SUMB_11_6_port);
   U56 : XOR2X1 port map( A => CARRYB_10_6_port, B => ab_11_6_port, Y => n34);
   U57 : XNOR2X1 port map( A => n508, B => n35, Y => SUMB_6_4_port);
   U58 : INVX1 port map( A => SUMB_5_5_port, Y => n35);
   U59 : XNOR2X1 port map( A => SUMB_8_4_port, B => n36, Y => SUMB_9_3_port);
   U60 : XNOR2X1 port map( A => CARRYB_8_3_port, B => ab_9_3_port, Y => n36);
   U61 : XOR2X1 port map( A => n37, B => n415, Y => SUMB_2_8_port);
   U62 : XOR2X1 port map( A => SUMB_1_9_port, B => ab_2_8_port, Y => n37);
   U63 : XOR2X1 port map( A => n38, B => ab_10_1_port, Y => n40);
   U64 : INVX1 port map( A => SUMB_9_2_port, Y => n38);
   U65 : XOR2X1 port map( A => n39, B => n40, Y => SUMB_10_1_port);
   U66 : INVX1 port map( A => n7, Y => n39);
   U67 : XOR2X1 port map( A => SUMB_6_10_port, B => n107, Y => n41);
   U68 : XNOR2X1 port map( A => n42, B => SUMB_3_11_port, Y => SUMB_4_10_port);
   U69 : XNOR2X1 port map( A => ab_4_10_port, B => CARRYB_3_10_port, Y => n42);
   U70 : XOR2X1 port map( A => n43, B => SUMB_8_9_port, Y => SUMB_9_8_port);
   U71 : XNOR2X1 port map( A => n248, B => CARRYB_8_8_port, Y => n43);
   U72 : NAND3X1 port map( A => n483, B => n482, C => n484, Y => n44);
   U73 : NAND3X1 port map( A => n865, B => n866, C => n867, Y => n45);
   U74 : INVX1 port map( A => SUMB_15_4_port, Y => n46);
   U75 : INVX1 port map( A => n46, Y => n47);
   U76 : BUFX4 port map( A => n1016, Y => n655);
   U77 : NAND3X1 port map( A => n561, B => n560, C => n562, Y => n48);
   U78 : NAND3X1 port map( A => n156, B => n155, C => n157, Y => n49);
   U79 : NAND3X1 port map( A => n939, B => n940, C => n941, Y => n50);
   U80 : NAND3X1 port map( A => n546, B => n545, C => n547, Y => n51);
   U81 : BUFX2 port map( A => CARRYB_9_0_port, Y => n52);
   U82 : BUFX2 port map( A => CARRYB_6_1_port, Y => n53);
   U83 : NAND3X1 port map( A => n856, B => n857, C => n858, Y => n54);
   U84 : NAND3X1 port map( A => n805, B => n806, C => n807, Y => n55);
   U85 : NAND3X1 port map( A => n574, B => n572, C => n573, Y => n56);
   U86 : NAND3X1 port map( A => n379, B => n378, C => n380, Y => n57);
   U87 : XNOR2X1 port map( A => CARRYB_7_6_port, B => n58, Y => n447);
   U88 : INVX8 port map( A => n104, Y => n58);
   U89 : INVX4 port map( A => n989, Y => n974);
   U90 : INVX4 port map( A => B(0), Y => n989);
   U91 : AND2X2 port map( A => ab_0_6_port, B => ab_1_5_port, Y => n59);
   U92 : NAND3X1 port map( A => n492, B => n493, C => n494, Y => n60);
   U93 : XOR2X1 port map( A => n61, B => n62, Y => SUMB_11_4_port);
   U94 : XNOR2X1 port map( A => n970, B => ab_11_4_port, Y => n61);
   U95 : XNOR2X1 port map( A => n220, B => n444, Y => n62);
   U96 : INVX2 port map( A => SUMB_12_2_port, Y => n400);
   U97 : INVX2 port map( A => SUMB_2_6_port, Y => n385);
   U98 : XOR2X1 port map( A => CARRYB_14_3_port, B => n63, Y => n595);
   U99 : INVX8 port map( A => ab_15_3_port, Y => n63);
   U100 : XNOR2X1 port map( A => n64, B => SUMB_10_6_port, Y => SUMB_11_5_port)
                           ;
   U101 : XNOR2X1 port map( A => CARRYB_10_5_port, B => ab_11_5_port, Y => n64)
                           ;
   U102 : INVX2 port map( A => SUMB_6_7_port, Y => n374);
   U103 : INVX2 port map( A => SUMB_12_4_port, Y => n221);
   U104 : XNOR2X1 port map( A => n65, B => SUMB_3_10_port, Y => SUMB_4_9_port);
   U105 : XNOR2X1 port map( A => n325, B => ab_4_9_port, Y => n65);
   U106 : INVX1 port map( A => n970, Y => n971);
   U107 : INVX2 port map( A => ab_8_8_port, Y => n280);
   U108 : INVX2 port map( A => ab_9_7_port, Y => n200);
   U109 : INVX2 port map( A => n414, Y => n178);
   U110 : INVX2 port map( A => ab_5_9_port, Y => n530);
   U111 : INVX2 port map( A => ab_3_12_port, Y => n150);
   U112 : INVX2 port map( A => ab_6_9_port, Y => n149);
   U113 : INVX2 port map( A => ab_10_5_port, Y => n130);
   U114 : INVX2 port map( A => ab_9_8_port, Y => n248);
   U115 : INVX2 port map( A => B(4), Y => n997);
   U116 : INVX2 port map( A => ab_13_5_port, Y => n201);
   U117 : INVX2 port map( A => ab_12_7_port, Y => n568);
   U118 : INVX2 port map( A => ab_5_8_port, Y => n362);
   U119 : INVX2 port map( A => ab_6_8_port, Y => n162);
   U120 : INVX2 port map( A => ab_4_6_port, Y => n317);
   U121 : INVX2 port map( A => ab_3_5_port, Y => n250);
   U122 : INVX2 port map( A => ab_2_15_port, Y => n243);
   U123 : INVX2 port map( A => ab_8_6_port, Y => n104);
   U124 : INVX2 port map( A => ab_5_10_port, Y => n279);
   U125 : INVX2 port map( A => ab_4_3_port, Y => n501);
   U126 : INVX2 port map( A => ab_8_4_port, Y => n175);
   U127 : INVX2 port map( A => ab_12_3_port, Y => n222);
   U128 : INVX2 port map( A => ab_6_10_port, Y => n247);
   U129 : INVX2 port map( A => ab_15_2_port, Y => n476);
   U130 : INVX1 port map( A => SUMB_6_14_port, Y => n296);
   U131 : INVX2 port map( A => ab_15_4_port, Y => n210);
   U132 : INVX2 port map( A => ab_12_1_port, Y => n804);
   U133 : INVX2 port map( A => CARRYB_15_6_port, Y => n294);
   U134 : INVX2 port map( A => B(11), Y => n1008);
   U135 : INVX4 port map( A => n1010, Y => n1011);
   U136 : INVX2 port map( A => B(14), Y => n1014);
   U137 : AND2X2 port map( A => SUMB_15_9_port, B => CARRYB_15_8_port, Y => n66
                           );
   U138 : AND2X2 port map( A => SUMB_15_10_port, B => CARRYB_15_9_port, Y => 
                           n67);
   U139 : AND2X2 port map( A => SUMB_15_11_port, B => CARRYB_15_10_port, Y => 
                           n68);
   U140 : AND2X2 port map( A => SUMB_15_12_port, B => CARRYB_15_11_port, Y => 
                           n69);
   U141 : AND2X2 port map( A => SUMB_15_13_port, B => CARRYB_15_12_port, Y => 
                           n70);
   U142 : AND2X2 port map( A => SUMB_15_14_port, B => CARRYB_15_13_port, Y => 
                           n71);
   U143 : AND2X2 port map( A => SUMB_15_15_port, B => CARRYB_15_14_port, Y => 
                           n72);
   U144 : INVX1 port map( A => CARRYB_3_1_port, Y => n988);
   U145 : INVX1 port map( A => CARRYB_6_13_port, Y => n368);
   U146 : AND2X2 port map( A => ab_1_7_port, B => ab_0_8_port, Y => n73);
   U147 : INVX2 port map( A => n959, Y => n979);
   U148 : INVX2 port map( A => B(10), Y => n1006);
   U149 : INVX2 port map( A => ab_13_3_port, Y => n477);
   U150 : XOR2X1 port map( A => n412, B => n74, Y => SUMB_8_1_port);
   U151 : XNOR2X1 port map( A => CARRYB_7_1_port, B => ab_8_1_port, Y => n74);
   U152 : BUFX2 port map( A => SUMB_4_4_port, Y => n75);
   U153 : BUFX2 port map( A => SUMB_13_2_port, Y => n76);
   U154 : BUFX2 port map( A => SUMB_4_11_port, Y => n77);
   U155 : BUFX2 port map( A => CARRYB_3_2_port, Y => n78);
   U156 : XOR2X1 port map( A => n143, B => n92, Y => n79);
   U157 : XNOR2X1 port map( A => n80, B => ab_0_14_port, Y => SUMB_1_13_port);
   U158 : NAND2X1 port map( A => n1018, B => n1013, Y => n80);
   U159 : BUFX2 port map( A => SUMB_8_2_port, Y => n81);
   U160 : NAND3X1 port map( A => n709, B => n710, C => n711, Y => n82);
   U161 : XNOR2X1 port map( A => n83, B => SUMB_12_6_port, Y => SUMB_13_5_port)
                           ;
   U162 : XOR2X1 port map( A => CARRYB_12_5_port, B => n201, Y => n83);
   U163 : XNOR2X1 port map( A => n84, B => CARRYB_5_9_port, Y => SUMB_6_9_port)
                           ;
   U164 : XOR2X1 port map( A => SUMB_5_10_port, B => n149, Y => n84);
   U165 : BUFX2 port map( A => CARRYB_7_0_port, Y => n85);
   U166 : BUFX2 port map( A => SUMB_7_1_port, Y => n86);
   U167 : NAND3X1 port map( A => n839, B => n838, C => n840, Y => n87);
   U168 : NAND3X1 port map( A => n781, B => n782, C => n783, Y => n88);
   U169 : XOR2X1 port map( A => n315, B => n442, Y => n89);
   U170 : INVX2 port map( A => SUMB_13_3_port, Y => n442);
   U171 : XOR2X1 port map( A => n90, B => SUMB_6_9_port, Y => SUMB_7_8_port);
   U172 : XOR2X1 port map( A => CARRYB_6_8_port, B => ab_7_8_port, Y => n90);
   U173 : XNOR2X1 port map( A => CARRYB_8_6_port, B => ab_9_6_port, Y => n148);
   U174 : BUFX2 port map( A => n864, Y => n91);
   U175 : BUFX2 port map( A => CARRYB_9_4_port, Y => n92);
   U176 : NAND3X1 port map( A => n868, B => n869, C => n870, Y => n93);
   U177 : NAND3X1 port map( A => n541, B => n542, C => n540, Y => n94);
   U178 : NAND3X1 port map( A => n659, B => n660, C => n661, Y => n95);
   U179 : NOR2X1 port map( A => n1012, B => n655, Y => n96);
   U180 : NAND3X1 port map( A => n827, B => n828, C => n829, Y => n97);
   U181 : BUFX2 port map( A => SUMB_2_5_port, Y => n98);
   U182 : XNOR2X1 port map( A => n99, B => n59, Y => SUMB_2_5_port);
   U183 : XNOR2X1 port map( A => SUMB_1_6_port, B => ab_2_5_port, Y => n99);
   U184 : XOR2X1 port map( A => n100, B => n385, Y => SUMB_3_5_port);
   U185 : XOR2X1 port map( A => CARRYB_2_5_port, B => n250, Y => n100);
   U186 : NAND2X1 port map( A => n765, B => n767, Y => n101);
   U187 : INVX2 port map( A => n101, Y => n102);
   U188 : INVX2 port map( A => CARRYB_15_4_port, Y => n293);
   U189 : XOR2X1 port map( A => n103, B => n158, Y => SUMB_5_5_port);
   U190 : XNOR2X1 port map( A => CARRYB_4_5_port, B => ab_5_5_port, Y => n103);
   U191 : XNOR2X1 port map( A => n105, B => SUMB_11_5_port, Y => SUMB_12_4_port
                           );
   U192 : XNOR2X1 port map( A => CARRYB_11_4_port, B => ab_12_4_port, Y => n105
                           );
   U193 : BUFX2 port map( A => SUMB_3_9_port, Y => n106);
   U194 : XOR2X1 port map( A => CARRYB_6_9_port, B => ab_7_9_port, Y => n107);
   U195 : XOR2X1 port map( A => SUMB_6_10_port, B => n107, Y => SUMB_7_9_port);
   U196 : NAND2X1 port map( A => SUMB_6_10_port, B => CARRYB_6_9_port, Y => 
                           n108);
   U197 : NAND2X1 port map( A => SUMB_6_10_port, B => ab_7_9_port, Y => n109);
   U198 : NAND2X1 port map( A => CARRYB_6_9_port, B => ab_7_9_port, Y => n110);
   U199 : NAND3X1 port map( A => n109, B => n108, C => n110, Y => 
                           CARRYB_7_9_port);
   U200 : NAND3X1 port map( A => n821, B => n822, C => n823, Y => n111);
   U201 : NAND3X1 port map( A => n818, B => n819, C => n820, Y => n112);
   U202 : XOR2X1 port map( A => ab_14_8_port, B => CARRYB_13_8_port, Y => n113)
                           ;
   U203 : XOR2X1 port map( A => n113, B => SUMB_13_9_port, Y => SUMB_14_8_port)
                           ;
   U204 : XOR2X1 port map( A => ab_15_7_port, B => CARRYB_14_7_port, Y => n114)
                           ;
   U205 : XOR2X1 port map( A => n114, B => SUMB_14_8_port, Y => SUMB_15_7_port)
                           ;
   U206 : NAND2X1 port map( A => ab_14_8_port, B => CARRYB_13_8_port, Y => n115
                           );
   U207 : NAND2X1 port map( A => ab_14_8_port, B => SUMB_13_9_port, Y => n116);
   U208 : NAND2X1 port map( A => CARRYB_13_8_port, B => SUMB_13_9_port, Y => 
                           n117);
   U209 : NAND3X1 port map( A => n115, B => n116, C => n117, Y => 
                           CARRYB_14_8_port);
   U210 : NAND2X1 port map( A => ab_15_7_port, B => CARRYB_14_7_port, Y => n118
                           );
   U211 : NAND2X1 port map( A => ab_15_7_port, B => SUMB_14_8_port, Y => n119);
   U212 : NAND2X1 port map( A => CARRYB_14_7_port, B => SUMB_14_8_port, Y => 
                           n120);
   U213 : NAND3X1 port map( A => n118, B => n119, C => n120, Y => 
                           CARRYB_15_7_port);
   U214 : XOR2X1 port map( A => SUMB_8_11_port, B => ab_9_10_port, Y => n121);
   U215 : XOR2X1 port map( A => n121, B => CARRYB_8_10_port, Y => 
                           SUMB_9_10_port);
   U216 : NAND2X1 port map( A => CARRYB_8_10_port, B => SUMB_8_11_port, Y => 
                           n122);
   U217 : NAND2X1 port map( A => CARRYB_8_10_port, B => ab_9_10_port, Y => n123
                           );
   U218 : NAND2X1 port map( A => SUMB_8_11_port, B => ab_9_10_port, Y => n124);
   U219 : NAND3X1 port map( A => n123, B => n122, C => n124, Y => 
                           CARRYB_9_10_port);
   U220 : XOR2X1 port map( A => CARRYB_12_8_port, B => ab_13_8_port, Y => n125)
                           ;
   U221 : XOR2X1 port map( A => SUMB_12_9_port, B => n125, Y => SUMB_13_8_port)
                           ;
   U222 : NAND2X1 port map( A => SUMB_12_9_port, B => CARRYB_12_8_port, Y => 
                           n126);
   U223 : NAND2X1 port map( A => SUMB_12_9_port, B => ab_13_8_port, Y => n127);
   U224 : NAND2X1 port map( A => CARRYB_12_8_port, B => ab_13_8_port, Y => n128
                           );
   U225 : NAND3X1 port map( A => n127, B => n126, C => n128, Y => 
                           CARRYB_13_8_port);
   U226 : NAND3X1 port map( A => n916, B => n915, C => n917, Y => n129);
   U227 : XNOR2X1 port map( A => CARRYB_9_5_port, B => n130, Y => n220);
   U228 : XOR2X1 port map( A => n131, B => n179, Y => SUMB_6_2_port);
   U229 : XOR2X1 port map( A => ab_6_2_port, B => n50, Y => n131);
   U230 : INVX4 port map( A => n991, Y => n980);
   U231 : INVX2 port map( A => n1016, Y => n401);
   U232 : INVX1 port map( A => n593, Y => n132);
   U233 : XNOR2X1 port map( A => n504, B => n254, Y => n133);
   U234 : NAND3X1 port map( A => n845, B => n847, C => n846, Y => n134);
   U235 : XNOR2X1 port map( A => n135, B => n136, Y => SUMB_12_2_port);
   U236 : XOR2X1 port map( A => CARRYB_11_2_port, B => ab_12_2_port, Y => n135)
                           ;
   U237 : INVX1 port map( A => SUMB_11_3_port, Y => n136);
   U238 : BUFX2 port map( A => SUMB_8_3_port, Y => n137);
   U239 : XNOR2X1 port map( A => n138, B => SUMB_7_4_port, Y => SUMB_8_3_port);
   U240 : XNOR2X1 port map( A => CARRYB_7_3_port, B => ab_8_3_port, Y => n138);
   U241 : AND2X2 port map( A => n1018, B => n1013, Y => n139);
   U242 : XOR2X1 port map( A => n140, B => n221, Y => SUMB_13_3_port);
   U243 : XOR2X1 port map( A => CARRYB_12_3_port, B => n477, Y => n140);
   U244 : XOR2X1 port map( A => n141, B => n142, Y => SUMB_7_3_port);
   U245 : XNOR2X1 port map( A => CARRYB_6_3_port, B => ab_7_3_port, Y => n141);
   U246 : INVX1 port map( A => SUMB_6_4_port, Y => n142);
   U247 : XOR2X1 port map( A => SUMB_9_5_port, B => ab_10_4_port, Y => n143);
   U248 : XOR2X1 port map( A => n143, B => n92, Y => SUMB_10_4_port);
   U249 : NAND2X1 port map( A => SUMB_9_5_port, B => CARRYB_9_4_port, Y => n144
                           );
   U250 : NAND2X1 port map( A => CARRYB_9_4_port, B => ab_10_4_port, Y => n145)
                           ;
   U251 : NAND2X1 port map( A => SUMB_9_5_port, B => ab_10_4_port, Y => n146);
   U252 : NAND3X1 port map( A => n145, B => n146, C => n144, Y => 
                           CARRYB_10_4_port);
   U253 : XOR2X1 port map( A => n148, B => n147, Y => SUMB_9_6_port);
   U254 : INVX2 port map( A => SUMB_8_7_port, Y => n147);
   U255 : INVX4 port map( A => n1006, Y => n1007);
   U256 : XOR2X1 port map( A => CARRYB_2_12_port, B => n150, Y => n151);
   U257 : XNOR2X1 port map( A => n151, B => SUMB_2_13_port, Y => SUMB_3_12_port
                           );
   U258 : INVX2 port map( A => CARRYB_7_9_port, Y => n289);
   U259 : XNOR2X1 port map( A => ab_1_10_port, B => n152, Y => SUMB_1_10_port);
   U260 : NAND2X1 port map( A => n1009, B => n401, Y => n152);
   U261 : XOR2X1 port map( A => CARRYB_4_7_port, B => ab_5_7_port, Y => n771);
   U262 : XNOR2X1 port map( A => n153, B => n465, Y => SUMB_2_9_port);
   U263 : XOR2X1 port map( A => ab_2_9_port, B => n760, Y => n153);
   U264 : NAND3X1 port map( A => n266, B => n265, C => n267, Y => n154);
   U265 : AND2X2 port map( A => CARRYB_15_3_port, B => n47, Y => n954);
   U266 : NAND2X1 port map( A => SUMB_8_4_port, B => n57, Y => n155);
   U267 : NAND2X1 port map( A => SUMB_8_4_port, B => ab_9_3_port, Y => n156);
   U268 : NAND2X1 port map( A => n57, B => ab_9_3_port, Y => n157);
   U269 : NAND3X1 port map( A => n156, B => n155, C => n157, Y => 
                           CARRYB_9_3_port);
   U270 : INVX2 port map( A => SUMB_4_6_port, Y => n158);
   U271 : NAND3X1 port map( A => n656, B => n657, C => n658, Y => n159);
   U272 : BUFX2 port map( A => n903, Y => n161);
   U273 : XOR2X1 port map( A => CARRYB_7_7_port, B => ab_8_7_port, Y => n575);
   U274 : XOR2X1 port map( A => CARRYB_5_8_port, B => n162, Y => n307);
   U275 : BUFX2 port map( A => n1009, Y => n163);
   U276 : INVX4 port map( A => n1008, Y => n1009);
   U277 : NAND3X1 port map( A => n311, B => n310, C => n312, Y => n164);
   U278 : NAND3X1 port map( A => n436, B => n437, C => n438, Y => n165);
   U279 : XNOR2X1 port map( A => n166, B => n167, Y => SUMB_6_6_port);
   U280 : XOR2X1 port map( A => SUMB_5_7_port, B => ab_6_6_port, Y => n166);
   U281 : INVX1 port map( A => CARRYB_5_6_port, Y => n167);
   U282 : XNOR2X1 port map( A => n883, B => n168, Y => SUMB_12_1_port);
   U283 : INVX2 port map( A => SUMB_11_2_port, Y => n168);
   U284 : XOR2X1 port map( A => CARRYB_6_10_port, B => ab_7_10_port, Y => n169)
                           ;
   U285 : XOR2X1 port map( A => SUMB_6_11_port, B => n169, Y => SUMB_7_10_port)
                           ;
   U286 : NAND2X1 port map( A => SUMB_6_11_port, B => n54, Y => n170);
   U287 : NAND2X1 port map( A => SUMB_6_11_port, B => ab_7_10_port, Y => n171);
   U288 : NAND2X1 port map( A => n54, B => ab_7_10_port, Y => n172);
   U289 : NAND3X1 port map( A => n171, B => n170, C => n172, Y => 
                           CARRYB_7_10_port);
   U290 : XNOR2X1 port map( A => n173, B => n240, Y => SUMB_4_6_port);
   U291 : XNOR2X1 port map( A => n841, B => n317, Y => n173);
   U292 : INVX1 port map( A => SUMB_3_6_port, Y => n174);
   U293 : XOR2X1 port map( A => CARRYB_7_4_port, B => n175, Y => n373);
   U294 : BUFX2 port map( A => SUMB_2_2_port, Y => n176);
   U295 : INVX2 port map( A => n182, Y => n183);
   U296 : XNOR2X1 port map( A => n177, B => SUMB_13_7_port, Y => SUMB_14_6_port
                           );
   U297 : XNOR2X1 port map( A => ab_14_6_port, B => CARRYB_13_6_port, Y => n177
                           );
   U298 : XOR2X1 port map( A => n460, B => n178, Y => n219);
   U299 : BUFX2 port map( A => SUMB_5_3_port, Y => n179);
   U300 : NAND3X1 port map( A => n936, B => n937, C => n938, Y => n180);
   U301 : INVX2 port map( A => ab_2_7_port, Y => n381);
   U302 : AND2X2 port map( A => n1009, B => n402, Y => n181);
   U303 : INVX1 port map( A => n802, Y => n182);
   U304 : XOR2X1 port map( A => ab_11_11_port, B => CARRYB_10_11_port, Y => 
                           n184);
   U305 : XOR2X1 port map( A => n184, B => SUMB_10_12_port, Y => 
                           SUMB_11_11_port);
   U306 : XOR2X1 port map( A => ab_12_10_port, B => CARRYB_11_10_port, Y => 
                           n185);
   U307 : XOR2X1 port map( A => n185, B => SUMB_11_11_port, Y => 
                           SUMB_12_10_port);
   U308 : NAND2X1 port map( A => ab_11_11_port, B => CARRYB_10_11_port, Y => 
                           n186);
   U309 : NAND2X1 port map( A => ab_11_11_port, B => SUMB_10_12_port, Y => n187
                           );
   U310 : NAND2X1 port map( A => CARRYB_10_11_port, B => SUMB_10_12_port, Y => 
                           n188);
   U311 : NAND3X1 port map( A => n186, B => n187, C => n188, Y => 
                           CARRYB_11_11_port);
   U312 : NAND2X1 port map( A => ab_12_10_port, B => CARRYB_11_10_port, Y => 
                           n189);
   U313 : NAND2X1 port map( A => ab_12_10_port, B => SUMB_11_11_port, Y => n190
                           );
   U314 : NAND2X1 port map( A => CARRYB_11_10_port, B => SUMB_11_11_port, Y => 
                           n191);
   U315 : NAND3X1 port map( A => n189, B => n190, C => n191, Y => 
                           CARRYB_12_10_port);
   U316 : XOR2X1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, Y => n192)
                           ;
   U317 : XOR2X1 port map( A => n192, B => SUMB_8_13_port, Y => SUMB_9_12_port)
                           ;
   U318 : XOR2X1 port map( A => ab_10_11_port, B => CARRYB_9_11_port, Y => n193
                           );
   U319 : XOR2X1 port map( A => n193, B => SUMB_9_12_port, Y => SUMB_10_11_port
                           );
   U320 : NAND2X1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, Y => n194
                           );
   U321 : NAND2X1 port map( A => ab_9_12_port, B => SUMB_8_13_port, Y => n195);
   U322 : NAND2X1 port map( A => CARRYB_8_12_port, B => SUMB_8_13_port, Y => 
                           n196);
   U323 : NAND3X1 port map( A => n194, B => n195, C => n196, Y => 
                           CARRYB_9_12_port);
   U324 : NAND2X1 port map( A => ab_10_11_port, B => CARRYB_9_11_port, Y => 
                           n197);
   U325 : NAND2X1 port map( A => ab_10_11_port, B => SUMB_9_12_port, Y => n198)
                           ;
   U326 : NAND2X1 port map( A => CARRYB_9_11_port, B => SUMB_9_12_port, Y => 
                           n199);
   U327 : NAND3X1 port map( A => n197, B => n198, C => n199, Y => 
                           CARRYB_10_11_port);
   U328 : XOR2X1 port map( A => CARRYB_3_11_port, B => ab_4_11_port, Y => n281)
                           ;
   U329 : XOR2X1 port map( A => CARRYB_8_7_port, B => n200, Y => n274);
   U330 : XOR2X1 port map( A => ab_11_10_port, B => CARRYB_10_10_port, Y => 
                           n202);
   U331 : XOR2X1 port map( A => n202, B => SUMB_10_11_port, Y => 
                           SUMB_11_10_port);
   U332 : XOR2X1 port map( A => ab_12_9_port, B => n216, Y => n203);
   U333 : XOR2X1 port map( A => n203, B => SUMB_11_10_port, Y => SUMB_12_9_port
                           );
   U334 : NAND2X1 port map( A => ab_11_10_port, B => CARRYB_10_10_port, Y => 
                           n204);
   U335 : NAND2X1 port map( A => ab_11_10_port, B => SUMB_10_11_port, Y => n205
                           );
   U336 : NAND2X1 port map( A => CARRYB_10_10_port, B => SUMB_10_11_port, Y => 
                           n206);
   U337 : NAND3X1 port map( A => n204, B => n205, C => n206, Y => 
                           CARRYB_11_10_port);
   U338 : NAND2X1 port map( A => ab_12_9_port, B => n216, Y => n207);
   U339 : NAND2X1 port map( A => ab_12_9_port, B => SUMB_11_10_port, Y => n208)
                           ;
   U340 : NAND2X1 port map( A => n216, B => SUMB_11_10_port, Y => n209);
   U341 : NAND3X1 port map( A => n207, B => n208, C => n209, Y => 
                           CARRYB_12_9_port);
   U342 : XNOR2X1 port map( A => CARRYB_14_4_port, B => n210, Y => n741);
   U343 : XOR2X1 port map( A => n211, B => n212, Y => SUMB_7_11_port);
   U344 : XNOR2X1 port map( A => ab_7_11_port, B => CARRYB_6_11_port, Y => n211
                           );
   U345 : INVX1 port map( A => SUMB_6_12_port, Y => n212);
   U346 : XNOR2X1 port map( A => n213, B => SUMB_8_12_port, Y => SUMB_9_11_port
                           );
   U347 : XNOR2X1 port map( A => ab_9_11_port, B => CARRYB_8_11_port, Y => n213
                           );
   U348 : NAND3X1 port map( A => n754, B => n755, C => n756, Y => n214);
   U349 : INVX2 port map( A => CARRYB_11_9_port, Y => n215);
   U350 : INVX4 port map( A => n215, Y => n216);
   U351 : AND2X1 port map( A => n132, B => n291, Y => n952);
   U352 : BUFX2 port map( A => n578, Y => n217);
   U353 : BUFX2 port map( A => n799, Y => n218);
   U354 : XNOR2X1 port map( A => n220, B => n444, Y => SUMB_10_5_port);
   U355 : XOR2X1 port map( A => SUMB_11_4_port, B => n222, Y => n229);
   U356 : XNOR2X1 port map( A => n481, B => n223, Y => SUMB_6_7_port);
   U357 : INVX1 port map( A => SUMB_5_8_port, Y => n223);
   U358 : BUFX2 port map( A => n800, Y => n224);
   U359 : XOR2X1 port map( A => CARRYB_9_6_port, B => ab_10_6_port, Y => n228);
   U360 : NAND2X1 port map( A => ab_14_2_port, B => n389, Y => n225);
   U361 : INVX2 port map( A => SUMB_6_6_port, Y => n308);
   U362 : XNOR2X1 port map( A => n226, B => SUMB_11_6_port, Y => SUMB_12_5_port
                           );
   U363 : XNOR2X1 port map( A => CARRYB_11_5_port, B => ab_12_5_port, Y => n226
                           );
   U364 : XOR2X1 port map( A => n227, B => n89, Y => SUMB_15_1_port);
   U365 : XOR2X1 port map( A => CARRYB_14_1_port, B => ab_15_1_port, Y => n227)
                           ;
   U366 : XOR2X1 port map( A => SUMB_9_7_port, B => n228, Y => SUMB_10_6_port);
   U367 : XNOR2X1 port map( A => n230, B => SUMB_13_6_port, Y => SUMB_14_5_port
                           );
   U368 : XNOR2X1 port map( A => n97, B => ab_14_5_port, Y => n230);
   U369 : NAND3X1 port map( A => n874, B => n872, C => n873, Y => n231);
   U370 : XOR2X1 port map( A => n232, B => n308, Y => SUMB_7_5_port);
   U371 : XNOR2X1 port map( A => CARRYB_6_5_port, B => ab_7_5_port, Y => n232);
   U372 : XNOR2X1 port map( A => n233, B => SUMB_9_11_port, Y => 
                           SUMB_10_10_port);
   U373 : XNOR2X1 port map( A => ab_10_10_port, B => CARRYB_9_10_port, Y => 
                           n233);
   U374 : BUFX2 port map( A => SUMB_15_5_port, Y => n234);
   U375 : NAND3X1 port map( A => n808, B => n809, C => n810, Y => n235);
   U376 : NAND3X1 port map( A => n816, B => n815, C => n817, Y => n236);
   U377 : NAND3X1 port map( A => n495, B => n497, C => n496, Y => n237);
   U378 : INVX2 port map( A => CARRYB_6_12_port, Y => n238);
   U379 : INVX4 port map( A => n238, Y => n239);
   U380 : XOR2X1 port map( A => n664, B => n459, Y => n240);
   U381 : INVX2 port map( A => CARRYB_5_13_port, Y => n241);
   U382 : INVX4 port map( A => n241, Y => n242);
   U383 : XOR2X1 port map( A => n244, B => n243, Y => SUMB_3_14_port);
   U384 : XNOR2X1 port map( A => ab_3_14_port, B => CARRYB_2_14_port, Y => n244
                           );
   U385 : NAND3X1 port map( A => n472, B => n471, C => n473, Y => n245);
   U386 : AND2X2 port map( A => n139, B => ab_0_14_port, Y => n246);
   U387 : XNOR2X1 port map( A => n247, B => n111, Y => n852);
   U388 : NAND3X1 port map( A => n911, B => n912, C => n913, Y => n249);
   U389 : NAND2X1 port map( A => SUMB_4_6_port, B => n56, Y => n251);
   U390 : NAND2X1 port map( A => SUMB_4_6_port, B => ab_5_5_port, Y => n252);
   U391 : NAND2X1 port map( A => n56, B => ab_5_5_port, Y => n253);
   U392 : NAND3X1 port map( A => n252, B => n251, C => n253, Y => 
                           CARRYB_5_5_port);
   U393 : NAND2X1 port map( A => n695, B => n694, Y => n254);
   U394 : NAND3X1 port map( A => n794, B => n793, C => n795, Y => n255);
   U395 : INVX1 port map( A => n404, Y => n256);
   U396 : INVX2 port map( A => SUMB_2_12_port, Y => n264);
   U397 : XOR2X1 port map( A => n51, B => ab_9_1_port, Y => n257);
   U398 : XOR2X1 port map( A => n81, B => n257, Y => SUMB_9_1_port);
   U399 : NAND2X1 port map( A => SUMB_8_2_port, B => CARRYB_8_1_port, Y => n258
                           );
   U400 : NAND2X1 port map( A => SUMB_8_2_port, B => ab_9_1_port, Y => n259);
   U401 : NAND2X1 port map( A => CARRYB_8_1_port, B => ab_9_1_port, Y => n260);
   U402 : NAND3X1 port map( A => n259, B => n258, C => n260, Y => 
                           CARRYB_9_1_port);
   U403 : NAND3X1 port map( A => n724, B => n722, C => n723, Y => n261);
   U404 : XOR2X1 port map( A => n53, B => n262, Y => SUMB_7_1_port);
   U405 : XOR2X1 port map( A => SUMB_6_2_port, B => ab_7_1_port, Y => n262);
   U406 : XNOR2X1 port map( A => n975, B => ab_3_4_port, Y => n624);
   U407 : XOR2X1 port map( A => n263, B => n264, Y => SUMB_3_11_port);
   U408 : XNOR2X1 port map( A => ab_3_11_port, B => n165, Y => n263);
   U409 : AND2X1 port map( A => n234, B => CARRYB_15_4_port, Y => n956);
   U410 : NAND2X1 port map( A => SUMB_10_6_port, B => n255, Y => n265);
   U411 : NAND2X1 port map( A => SUMB_10_6_port, B => ab_11_5_port, Y => n266);
   U412 : NAND2X1 port map( A => n255, B => ab_11_5_port, Y => n267);
   U413 : NAND3X1 port map( A => n266, B => n265, C => n267, Y => 
                           CARRYB_11_5_port);
   U414 : NAND3X1 port map( A => n813, B => n812, C => n814, Y => n268);
   U415 : XNOR2X1 port map( A => n269, B => SUMB_5_6_port, Y => SUMB_6_5_port);
   U416 : XOR2X1 port map( A => n662, B => ab_6_5_port, Y => n269);
   U417 : NAND3X1 port map( A => n679, B => n681, C => n680, Y => n270);
   U418 : NAND3X1 port map( A => n712, B => n713, C => n714, Y => n271);
   U419 : NAND3X1 port map( A => n778, B => n779, C => n780, Y => n272);
   U420 : NAND3X1 port map( A => n706, B => n707, C => n708, Y => n273);
   U421 : XNOR2X1 port map( A => n274, B => n6, Y => SUMB_9_7_port);
   U422 : NAND2X1 port map( A => SUMB_11_4_port, B => CARRYB_11_3_port, Y => 
                           n275);
   U423 : NAND2X1 port map( A => CARRYB_11_3_port, B => ab_12_3_port, Y => n276
                           );
   U424 : NAND2X1 port map( A => SUMB_11_4_port, B => ab_12_3_port, Y => n277);
   U425 : NAND3X1 port map( A => n276, B => n275, C => n277, Y => 
                           CARRYB_12_3_port);
   U426 : NAND3X1 port map( A => n419, B => n421, C => n420, Y => n278);
   U427 : XOR2X1 port map( A => SUMB_4_11_port, B => n279, Y => n803);
   U428 : XOR2X1 port map( A => CARRYB_7_8_port, B => n280, Y => n282);
   U429 : XOR2X1 port map( A => n281, B => SUMB_3_12_port, Y => SUMB_4_11_port)
                           ;
   U430 : XNOR2X1 port map( A => n282, B => n41, Y => SUMB_8_8_port);
   U431 : XNOR2X1 port map( A => n283, B => SUMB_4_9_port, Y => SUMB_5_8_port);
   U432 : XOR2X1 port map( A => CARRYB_4_8_port, B => n362, Y => n283);
   U433 : NAND3X1 port map( A => n787, B => n788, C => n789, Y => n284);
   U434 : INVX2 port map( A => SUMB_9_6_port, Y => n444);
   U435 : INVX2 port map( A => CARRYB_5_12_port, Y => n285);
   U436 : INVX4 port map( A => n285, Y => n286);
   U437 : XOR2X1 port map( A => n287, B => n106, Y => SUMB_4_8_port);
   U438 : XOR2X1 port map( A => CARRYB_3_8_port, B => ab_4_8_port, Y => n287);
   U439 : XOR2X1 port map( A => n288, B => SUMB_10_8_port, Y => SUMB_11_7_port)
                           ;
   U440 : XOR2X1 port map( A => CARRYB_10_7_port, B => ab_11_7_port, Y => n288)
                           ;
   U441 : XNOR2X1 port map( A => n290, B => n289, Y => SUMB_8_9_port);
   U442 : XOR2X1 port map( A => SUMB_7_10_port, B => ab_8_9_port, Y => n290);
   U443 : BUFX2 port map( A => SUMB_15_3_port, Y => n291);
   U444 : INVX1 port map( A => CARRYB_2_9_port, Y => n875);
   U445 : INVX1 port map( A => n875, Y => n876);
   U446 : XNOR2X1 port map( A => n292, B => SUMB_12_7_port, Y => SUMB_13_6_port
                           );
   U447 : XNOR2X1 port map( A => CARRYB_12_6_port, B => ab_13_6_port, Y => n292
                           );
   U448 : XNOR2X1 port map( A => SUMB_15_5_port, B => n293, Y => A1_18_port);
   U449 : XNOR2X1 port map( A => ab_7_13_port, B => n368, Y => n629);
   U450 : XNOR2X1 port map( A => SUMB_15_7_port, B => n294, Y => A1_20_port);
   U451 : XNOR2X1 port map( A => SUMB_3_13_port, B => n295, Y => SUMB_4_12_port
                           );
   U452 : XNOR2X1 port map( A => CARRYB_3_12_port, B => ab_4_12_port, Y => n295
                           );
   U453 : XNOR2X1 port map( A => n629, B => n296, Y => SUMB_7_13_port);
   U454 : NAND2X1 port map( A => SUMB_4_7_port, B => n284, Y => n297);
   U455 : NAND2X1 port map( A => SUMB_4_7_port, B => ab_5_6_port, Y => n298);
   U456 : NAND2X1 port map( A => n284, B => ab_5_6_port, Y => n299);
   U457 : NAND3X1 port map( A => n298, B => n297, C => n299, Y => 
                           CARRYB_5_6_port);
   U458 : NAND3X1 port map( A => n416, B => n417, C => n12, Y => n300);
   U459 : NAND3X1 port map( A => n791, B => n792, C => n790, Y => n301);
   U460 : XOR2X1 port map( A => n302, B => SUMB_14_1_port, Y => SUMB_15_0_port)
                           ;
   U461 : NAND2X1 port map( A => n231, B => SUMB_14_1_port, Y => n303);
   U462 : NAND2X1 port map( A => SUMB_14_1_port, B => ab_15_0_port, Y => n304);
   U463 : NAND2X1 port map( A => n231, B => ab_15_0_port, Y => n305);
   U464 : NAND3X1 port map( A => n304, B => n303, C => n305, Y => 
                           CARRYB_15_0_port);
   U465 : XNOR2X1 port map( A => n306, B => SUMB_14_6_port, Y => SUMB_15_5_port
                           );
   U466 : XNOR2X1 port map( A => CARRYB_14_5_port, B => ab_15_5_port, Y => n306
                           );
   U467 : XNOR2X1 port map( A => n307, B => SUMB_5_9_port, Y => SUMB_6_8_port);
   U468 : XNOR2X1 port map( A => n372, B => SUMB_13_5_port, Y => SUMB_14_4_port
                           );
   U469 : XOR2X1 port map( A => CARRYB_9_3_port, B => ab_10_3_port, Y => n314);
   U470 : XOR2X1 port map( A => SUMB_3_3_port, B => ab_4_2_port, Y => n309);
   U471 : XOR2X1 port map( A => n309, B => n78, Y => SUMB_4_2_port);
   U472 : NAND2X1 port map( A => CARRYB_3_2_port, B => SUMB_3_3_port, Y => n310
                           );
   U473 : NAND2X1 port map( A => CARRYB_3_2_port, B => ab_4_2_port, Y => n311);
   U474 : NAND2X1 port map( A => SUMB_3_3_port, B => ab_4_2_port, Y => n312);
   U475 : NAND3X1 port map( A => n311, B => n310, C => n312, Y => 
                           CARRYB_4_2_port);
   U476 : BUFX2 port map( A => CARRYB_11_0_port, Y => n313);
   U477 : XNOR2X1 port map( A => n314, B => n425, Y => SUMB_10_3_port);
   U478 : XOR2X1 port map( A => n315, B => n442, Y => SUMB_14_2_port);
   U479 : XNOR2X1 port map( A => n316, B => n79, Y => SUMB_11_3_port);
   U480 : XNOR2X1 port map( A => CARRYB_10_3_port, B => ab_11_3_port, Y => n316
                           );
   U481 : NAND3X1 port map( A => n583, B => n584, C => n585, Y => n318);
   U482 : XOR2X1 port map( A => CARRYB_2_6_port, B => n319, Y => n503);
   U483 : NAND2X1 port map( A => n1022, B => n969, Y => n319);
   U484 : NAND2X1 port map( A => ab_12_1_port, B => n982, Y => n320);
   U485 : BUFX2 port map( A => SUMB_4_3_port, Y => n321);
   U486 : BUFX2 port map( A => CARRYB_7_2_port, Y => n322);
   U487 : XOR2X1 port map( A => n503, B => n323, Y => SUMB_3_6_port);
   U488 : INVX2 port map( A => n1002, Y => n905);
   U489 : BUFX2 port map( A => n688, Y => n324);
   U490 : NAND3X1 port map( A => n599, B => n598, C => n597, Y => n325);
   U491 : XOR2X1 port map( A => CARRYB_14_6_port, B => ab_15_6_port, Y => n326)
                           ;
   U492 : XOR2X1 port map( A => SUMB_14_7_port, B => n326, Y => SUMB_15_6_port)
                           ;
   U493 : NAND2X1 port map( A => SUMB_14_7_port, B => n11, Y => n327);
   U494 : NAND2X1 port map( A => SUMB_14_7_port, B => ab_15_6_port, Y => n328);
   U495 : NAND2X1 port map( A => n11, B => ab_15_6_port, Y => n329);
   U496 : NAND3X1 port map( A => n328, B => n327, C => n329, Y => 
                           CARRYB_15_6_port);
   U497 : XOR2X1 port map( A => CARRYB_13_7_port, B => ab_14_7_port, Y => n330)
                           ;
   U498 : XOR2X1 port map( A => SUMB_13_8_port, B => n330, Y => SUMB_14_7_port)
                           ;
   U499 : NAND2X1 port map( A => SUMB_13_8_port, B => CARRYB_13_7_port, Y => 
                           n331);
   U500 : NAND2X1 port map( A => SUMB_13_8_port, B => ab_14_7_port, Y => n332);
   U501 : NAND2X1 port map( A => CARRYB_13_7_port, B => ab_14_7_port, Y => n333
                           );
   U502 : NAND3X1 port map( A => n332, B => n331, C => n333, Y => 
                           CARRYB_14_7_port);
   U503 : INVX2 port map( A => CARRYB_6_7_port, Y => n404);
   U504 : NAND3X1 port map( A => n925, B => n926, C => n927, Y => n334);
   U505 : NAND2X1 port map( A => ab_14_6_port, B => n60, Y => n335);
   U506 : NAND2X1 port map( A => ab_14_6_port, B => SUMB_13_7_port, Y => n336);
   U507 : NAND2X1 port map( A => n60, B => SUMB_13_7_port, Y => n337);
   U508 : NAND3X1 port map( A => n335, B => n336, C => n337, Y => 
                           CARRYB_14_6_port);
   U509 : NAND2X1 port map( A => ab_15_5_port, B => n237, Y => n338);
   U510 : NAND2X1 port map( A => SUMB_14_6_port, B => ab_15_5_port, Y => n339);
   U511 : NAND2X1 port map( A => n237, B => n22, Y => n340);
   U512 : NAND3X1 port map( A => n338, B => n339, C => n340, Y => 
                           CARRYB_15_5_port);
   U513 : NAND2X1 port map( A => n643, B => n342, Y => n343);
   U514 : NAND2X1 port map( A => n341, B => SUMB_12_8_port, Y => n344);
   U515 : NAND2X1 port map( A => n343, B => n344, Y => SUMB_13_7_port);
   U516 : INVX1 port map( A => n643, Y => n341);
   U517 : INVX1 port map( A => SUMB_12_8_port, Y => n342);
   U518 : NAND3X1 port map( A => n853, B => n854, C => n855, Y => n345);
   U519 : NAND3X1 port map( A => n908, B => n909, C => n910, Y => n346);
   U520 : INVX2 port map( A => SUMB_9_3_port, Y => n347);
   U521 : XOR2X1 port map( A => ab_2_2_port, B => n960, Y => n348);
   U522 : XOR2X1 port map( A => n348, B => SUMB_1_3_port, Y => SUMB_2_2_port);
   U523 : XOR2X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, Y => n349);
   U524 : XOR2X1 port map( A => n349, B => n176, Y => SUMB_3_1_port);
   U525 : NAND2X1 port map( A => ab_2_2_port, B => n960, Y => n350);
   U526 : NAND2X1 port map( A => ab_2_2_port, B => SUMB_1_3_port, Y => n351);
   U527 : NAND2X1 port map( A => n960, B => SUMB_1_3_port, Y => n352);
   U528 : NAND3X1 port map( A => n350, B => n351, C => n352, Y => 
                           CARRYB_2_2_port);
   U529 : NAND2X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, Y => n353);
   U530 : NAND2X1 port map( A => ab_3_1_port, B => SUMB_2_2_port, Y => n354);
   U531 : NAND2X1 port map( A => CARRYB_2_1_port, B => SUMB_2_2_port, Y => n355
                           );
   U532 : NAND3X1 port map( A => n353, B => n354, C => n355, Y => 
                           CARRYB_3_1_port);
   U533 : XOR2X1 port map( A => SUMB_10_1_port, B => ab_11_0_port, Y => n356);
   U534 : XOR2X1 port map( A => n967, B => n356, Y => A1_9_port);
   U535 : NAND2X1 port map( A => n967, B => SUMB_10_1_port, Y => n357);
   U536 : NAND2X1 port map( A => n967, B => ab_11_0_port, Y => n358);
   U537 : NAND2X1 port map( A => SUMB_10_1_port, B => ab_11_0_port, Y => n359);
   U538 : NAND3X1 port map( A => n358, B => n357, C => n359, Y => 
                           CARRYB_11_0_port);
   U539 : BUFX2 port map( A => SUMB_4_1_port, Y => n360);
   U540 : XNOR2X1 port map( A => n361, B => SUMB_10_9_port, Y => SUMB_11_8_port
                           );
   U541 : XNOR2X1 port map( A => ab_11_8_port, B => CARRYB_10_8_port, Y => n361
                           );
   U542 : XNOR2X1 port map( A => n934, B => n363, Y => SUMB_4_3_port);
   U543 : INVX2 port map( A => SUMB_3_4_port, Y => n363);
   U544 : XOR2X1 port map( A => n364, B => n365, Y => SUMB_11_2_port);
   U545 : XNOR2X1 port map( A => ab_11_2_port, B => CARRYB_10_2_port, Y => n364
                           );
   U546 : INVX1 port map( A => SUMB_10_3_port, Y => n365);
   U547 : INVX2 port map( A => CARRYB_4_13_port, Y => n366);
   U548 : INVX4 port map( A => n366, Y => n367);
   U549 : NAND3X1 port map( A => n796, B => n797, C => n798, Y => n369);
   U550 : XOR2X1 port map( A => n28, B => n370, Y => SUMB_13_2_port);
   U551 : XOR2X1 port map( A => CARRYB_12_2_port, B => ab_13_2_port, Y => n370)
                           ;
   U552 : XOR2X1 port map( A => n606, B => n371, Y => SUMB_8_5_port);
   U553 : INVX1 port map( A => SUMB_7_6_port, Y => n371);
   U554 : XNOR2X1 port map( A => CARRYB_13_4_port, B => ab_14_4_port, Y => n372
                           );
   U555 : XOR2X1 port map( A => n737, B => n375, Y => SUMB_4_7_port);
   U556 : INVX1 port map( A => SUMB_3_8_port, Y => n375);
   U557 : XNOR2X1 port map( A => ab_2_13_port, B => n966, Y => n914);
   U558 : INVX2 port map( A => n570, Y => n571);
   U559 : NAND3X1 port map( A => n791, B => n792, C => n790, Y => n376);
   U560 : NAND3X1 port map( A => n894, B => n896, C => n895, Y => n377);
   U561 : NAND2X1 port map( A => SUMB_7_4_port, B => CARRYB_7_3_port, Y => n378
                           );
   U562 : NAND2X1 port map( A => SUMB_7_4_port, B => ab_8_3_port, Y => n379);
   U563 : NAND2X1 port map( A => CARRYB_7_3_port, B => ab_8_3_port, Y => n380);
   U564 : NAND3X1 port map( A => n379, B => n378, C => n380, Y => 
                           CARRYB_8_3_port);
   U565 : XOR2X1 port map( A => n906, B => n381, Y => n468);
   U566 : NAND2X1 port map( A => n59, B => SUMB_1_6_port, Y => n382);
   U567 : NAND2X1 port map( A => n59, B => ab_2_5_port, Y => n383);
   U568 : NAND2X1 port map( A => SUMB_1_6_port, B => ab_2_5_port, Y => n384);
   U569 : NAND3X1 port map( A => n383, B => n382, C => n384, Y => 
                           CARRYB_2_5_port);
   U570 : AND2X2 port map( A => B(7), B => A(2), Y => ab_2_7_port);
   U571 : NAND3X1 port map( A => n889, B => n890, C => n888, Y => n386);
   U572 : NAND3X1 port map( A => n945, B => n946, C => n947, Y => n387);
   U573 : NAND3X1 port map( A => n553, B => n551, C => n552, Y => n388);
   U574 : NAND3X1 port map( A => n920, B => n921, C => n919, Y => n389);
   U575 : NAND3X1 port map( A => n893, B => n892, C => n891, Y => n390);
   U576 : NAND3X1 port map( A => n801, B => n218, C => n224, Y => n391);
   U577 : NAND3X1 port map( A => n687, B => n324, C => n689, Y => n392);
   U578 : NAND3X1 port map( A => n862, B => n91, C => n863, Y => n393);
   U579 : NAND3X1 port map( A => n901, B => n902, C => n161, Y => n394);
   U580 : NAND3X1 port map( A => n842, B => n843, C => n844, Y => n395);
   U581 : NAND3X1 port map( A => n556, B => n554, C => n555, Y => n396);
   U582 : NAND3X1 port map( A => n922, B => n923, C => n924, Y => n397);
   U583 : NAND3X1 port map( A => n768, B => n769, C => n770, Y => n398);
   U584 : BUFX2 port map( A => n577, Y => n399);
   U585 : XNOR2X1 port map( A => n705, B => ab_7_2_port, Y => n449);
   U586 : XNOR2X1 port map( A => n837, B => n400, Y => SUMB_13_1_port);
   U587 : INVX2 port map( A => n1016, Y => n402);
   U588 : INVX2 port map( A => B(12), Y => n1010);
   U589 : XOR2X1 port map( A => n664, B => n459, Y => SUMB_3_7_port);
   U590 : NAND2X1 port map( A => ab_7_7_port, B => n404, Y => n405);
   U591 : NAND2X1 port map( A => n403, B => n44, Y => n406);
   U592 : NAND2X1 port map( A => n405, B => n406, Y => n897);
   U593 : INVX1 port map( A => ab_7_7_port, Y => n403);
   U594 : NAND3X1 port map( A => n587, B => n588, C => n589, Y => n407);
   U595 : XOR2X1 port map( A => SUMB_9_1_port, B => ab_10_0_port, Y => n408);
   U596 : XOR2X1 port map( A => n52, B => n408, Y => A1_8_port);
   U597 : NAND2X1 port map( A => CARRYB_9_0_port, B => SUMB_9_1_port, Y => n409
                           );
   U598 : NAND2X1 port map( A => CARRYB_9_0_port, B => ab_10_0_port, Y => n410)
                           ;
   U599 : NAND2X1 port map( A => SUMB_9_1_port, B => ab_10_0_port, Y => n411);
   U600 : NAND3X1 port map( A => n410, B => n409, C => n411, Y => 
                           CARRYB_10_0_port);
   U601 : INVX1 port map( A => SUMB_7_2_port, Y => n412);
   U602 : INVX8 port map( A => n1017, Y => n1018);
   U603 : XNOR2X1 port map( A => n413, B => SUMB_2_4_port, Y => SUMB_3_3_port);
   U604 : XOR2X1 port map( A => n983, B => ab_3_3_port, Y => n413);
   U605 : INVX2 port map( A => n478, Y => n414);
   U606 : NOR2X1 port map( A => n1017, B => n1008, Y => ab_1_11_port);
   U607 : XNOR2X1 port map( A => n460, B => n414, Y => SUMB_2_10_port);
   U608 : AND2X2 port map( A => ab_1_8_port, B => ab_0_9_port, Y => n415);
   U609 : NAND2X1 port map( A => SUMB_5_7_port, B => ab_6_6_port, Y => n416);
   U610 : NAND2X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, Y => n417);
   U611 : NAND2X1 port map( A => SUMB_5_7_port, B => CARRYB_5_6_port, Y => n418
                           );
   U612 : NAND3X1 port map( A => n417, B => n416, C => n418, Y => 
                           CARRYB_6_6_port);
   U613 : NAND2X1 port map( A => ab_7_5_port, B => n334, Y => n419);
   U614 : NAND2X1 port map( A => SUMB_6_6_port, B => ab_7_5_port, Y => n420);
   U615 : NAND2X1 port map( A => SUMB_6_6_port, B => n334, Y => n421);
   U616 : NAND3X1 port map( A => n421, B => n420, C => n419, Y => 
                           CARRYB_7_5_port);
   U617 : XNOR2X1 port map( A => n422, B => SUMB_2_9_port, Y => SUMB_3_8_port);
   U618 : XNOR2X1 port map( A => n376, B => n538, Y => n422);
   U619 : XOR2X1 port map( A => n424, B => SUMB_6_5_port, Y => SUMB_7_4_port);
   U620 : XOR2X1 port map( A => CARRYB_6_4_port, B => ab_7_4_port, Y => n424);
   U621 : INVX1 port map( A => SUMB_9_4_port, Y => n425);
   U622 : XOR2X1 port map( A => CARRYB_13_1_port, B => ab_14_1_port, Y => n918)
                           ;
   U623 : XOR2X1 port map( A => n48, B => ab_3_9_port, Y => n596);
   U624 : XOR2X1 port map( A => CARRYB_2_13_port, B => ab_3_13_port, Y => n426)
                           ;
   U625 : XOR2X1 port map( A => SUMB_2_14_port, B => n426, Y => SUMB_3_13_port)
                           ;
   U626 : NAND2X1 port map( A => SUMB_2_14_port, B => n129, Y => n427);
   U627 : NAND2X1 port map( A => SUMB_2_14_port, B => ab_3_13_port, Y => n428);
   U628 : NAND2X1 port map( A => n129, B => ab_3_13_port, Y => n429);
   U629 : NAND3X1 port map( A => n428, B => n427, C => n429, Y => 
                           CARRYB_3_13_port);
   U630 : XOR2X1 port map( A => ab_1_15_port, B => ab_2_14_port, Y => n430);
   U631 : XOR2X1 port map( A => n430, B => n30, Y => SUMB_2_14_port);
   U632 : NAND2X1 port map( A => n961, B => ab_1_15_port, Y => n431);
   U633 : NAND2X1 port map( A => n961, B => ab_2_14_port, Y => n432);
   U634 : NAND2X1 port map( A => ab_1_15_port, B => ab_2_14_port, Y => n433);
   U635 : NAND3X1 port map( A => n432, B => n431, C => n433, Y => 
                           CARRYB_2_14_port);
   U636 : XOR2X1 port map( A => ab_2_11_port, B => n506, Y => n434);
   U637 : XOR2X1 port map( A => n434, B => SUMB_1_12_port, Y => SUMB_2_11_port)
                           ;
   U638 : XOR2X1 port map( A => ab_3_10_port, B => CARRYB_2_10_port, Y => n435)
                           ;
   U639 : XOR2X1 port map( A => n435, B => SUMB_2_11_port, Y => SUMB_3_10_port)
                           ;
   U640 : NAND2X1 port map( A => ab_2_11_port, B => n506, Y => n436);
   U641 : NAND2X1 port map( A => ab_2_11_port, B => SUMB_1_12_port, Y => n437);
   U642 : NAND2X1 port map( A => n506, B => SUMB_1_12_port, Y => n438);
   U643 : NAND3X1 port map( A => n436, B => n437, C => n438, Y => 
                           CARRYB_2_11_port);
   U644 : NAND2X1 port map( A => ab_3_10_port, B => CARRYB_2_10_port, Y => n439
                           );
   U645 : NAND2X1 port map( A => ab_3_10_port, B => SUMB_2_11_port, Y => n440);
   U646 : NAND2X1 port map( A => CARRYB_2_10_port, B => SUMB_2_11_port, Y => 
                           n441);
   U647 : NAND3X1 port map( A => n439, B => n440, C => n441, Y => 
                           CARRYB_3_10_port);
   U648 : NAND3X1 port map( A => n775, B => n777, C => n776, Y => n443);
   U649 : INVX2 port map( A => SUMB_7_7_port, Y => n448);
   U650 : BUFX2 port map( A => SUMB_1_5_port, Y => n445);
   U651 : BUFX2 port map( A => CARRYB_3_6_port, Y => n446);
   U652 : XOR2X1 port map( A => n447, B => n448, Y => SUMB_8_6_port);
   U653 : XOR2X1 port map( A => SUMB_6_3_port, B => n449, Y => SUMB_7_2_port);
   U654 : NAND2X1 port map( A => SUMB_6_3_port, B => CARRYB_6_2_port, Y => n450
                           );
   U655 : NAND2X1 port map( A => SUMB_6_3_port, B => ab_7_2_port, Y => n451);
   U656 : NAND2X1 port map( A => CARRYB_6_2_port, B => ab_7_2_port, Y => n452);
   U657 : NAND3X1 port map( A => n451, B => n450, C => n452, Y => 
                           CARRYB_7_2_port);
   U658 : XOR2X1 port map( A => CARRYB_8_2_port, B => ab_9_2_port, Y => n453);
   U659 : XOR2X1 port map( A => n453, B => n137, Y => SUMB_9_2_port);
   U660 : NAND2X1 port map( A => SUMB_8_3_port, B => n458, Y => n454);
   U661 : NAND2X1 port map( A => SUMB_8_3_port, B => ab_9_2_port, Y => n455);
   U662 : NAND2X1 port map( A => n458, B => ab_9_2_port, Y => n456);
   U663 : NAND3X1 port map( A => n455, B => n454, C => n456, Y => 
                           CARRYB_9_2_port);
   U664 : NAND3X1 port map( A => n532, B => n533, C => n534, Y => n457);
   U665 : NAND3X1 port map( A => n565, B => n564, C => n566, Y => n458);
   U666 : INVX2 port map( A => SUMB_2_8_port, Y => n459);
   U667 : XOR2X1 port map( A => SUMB_1_11_port, B => ab_2_10_port, Y => n460);
   U668 : NAND2X1 port map( A => SUMB_1_11_port, B => n478, Y => n461);
   U669 : NAND2X1 port map( A => n478, B => ab_2_10_port, Y => n462);
   U670 : NAND2X1 port map( A => SUMB_1_11_port, B => ab_2_10_port, Y => n463);
   U671 : NAND3X1 port map( A => n462, B => n461, C => n463, Y => 
                           CARRYB_2_10_port);
   U672 : XNOR2X1 port map( A => n395, B => ab_13_4_port, Y => n464);
   U673 : INVX1 port map( A => SUMB_1_10_port, Y => n465);
   U674 : NAND3X1 port map( A => n898, B => n899, C => n900, Y => n466);
   U675 : NAND3X1 port map( A => n579, B => n581, C => n580, Y => n467);
   U676 : XNOR2X1 port map( A => n468, B => SUMB_1_8_port, Y => SUMB_2_7_port);
   U677 : BUFX2 port map( A => SUMB_4_5_port, Y => n469);
   U678 : XOR2X1 port map( A => SUMB_1_7_port, B => ab_2_6_port, Y => n470);
   U679 : XOR2X1 port map( A => n470, B => n904, Y => SUMB_2_6_port);
   U680 : NAND2X1 port map( A => SUMB_1_7_port, B => n904, Y => n471);
   U681 : NAND2X1 port map( A => n904, B => ab_2_6_port, Y => n472);
   U682 : NAND2X1 port map( A => SUMB_1_7_port, B => ab_2_6_port, Y => n473);
   U683 : NAND3X1 port map( A => n472, B => n471, C => n473, Y => 
                           CARRYB_2_6_port);
   U684 : NAND3X1 port map( A => n225, B => n486, C => n487, Y => n474);
   U685 : NAND3X1 port map( A => n784, B => n785, C => n786, Y => n475);
   U686 : XNOR2X1 port map( A => CARRYB_14_2_port, B => n476, Y => n686);
   U687 : AND2X2 port map( A => n181, B => ab_1_10_port, Y => n478);
   U688 : NAND3X1 port map( A => n590, B => n591, C => n592, Y => n479);
   U689 : NAND3X1 port map( A => n576, B => n399, C => n217, Y => n480);
   U690 : XOR2X1 port map( A => n443, B => ab_6_7_port, Y => n481);
   U691 : NAND2X1 port map( A => SUMB_5_8_port, B => CARRYB_5_7_port, Y => n482
                           );
   U692 : NAND2X1 port map( A => SUMB_5_8_port, B => ab_6_7_port, Y => n483);
   U693 : NAND2X1 port map( A => CARRYB_5_7_port, B => ab_6_7_port, Y => n484);
   U694 : NAND3X1 port map( A => n483, B => n482, C => n484, Y => 
                           CARRYB_6_7_port);
   U695 : NAND2X1 port map( A => ab_14_2_port, B => n389, Y => n485);
   U696 : NAND2X1 port map( A => SUMB_13_3_port, B => ab_14_2_port, Y => n486);
   U697 : NAND2X1 port map( A => SUMB_13_3_port, B => n389, Y => n487);
   U698 : NAND3X1 port map( A => n485, B => n486, C => n487, Y => 
                           CARRYB_14_2_port);
   U699 : NAND2X1 port map( A => ab_15_1_port, B => n397, Y => n488);
   U700 : NAND2X1 port map( A => SUMB_14_2_port, B => ab_15_1_port, Y => n489);
   U701 : NAND2X1 port map( A => SUMB_14_2_port, B => n397, Y => n490);
   U702 : NAND3X1 port map( A => n488, B => n490, C => n489, Y => 
                           CARRYB_15_1_port);
   U703 : INVX4 port map( A => n997, Y => n977);
   U704 : INVX4 port map( A => A(3), Y => n1021);
   U705 : XNOR2X1 port map( A => n491, B => n75, Y => SUMB_5_3_port);
   U706 : XNOR2X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, Y => n491);
   U707 : NAND2X1 port map( A => ab_13_6_port, B => CARRYB_12_6_port, Y => n492
                           );
   U708 : NAND2X1 port map( A => SUMB_12_7_port, B => ab_13_6_port, Y => n493);
   U709 : NAND2X1 port map( A => CARRYB_12_6_port, B => SUMB_12_7_port, Y => 
                           n494);
   U710 : NAND3X1 port map( A => n492, B => n493, C => n494, Y => 
                           CARRYB_13_6_port);
   U711 : NAND2X1 port map( A => ab_14_5_port, B => n97, Y => n495);
   U712 : NAND2X1 port map( A => SUMB_13_6_port, B => ab_14_5_port, Y => n496);
   U713 : NAND2X1 port map( A => n97, B => SUMB_13_6_port, Y => n497);
   U714 : NAND3X1 port map( A => n495, B => n496, C => n497, Y => 
                           CARRYB_14_5_port);
   U715 : NAND2X1 port map( A => SUMB_10_8_port, B => n235, Y => n498);
   U716 : NAND2X1 port map( A => SUMB_10_8_port, B => ab_11_7_port, Y => n499);
   U717 : NAND2X1 port map( A => n235, B => ab_11_7_port, Y => n500);
   U718 : NAND3X1 port map( A => n499, B => n498, C => n500, Y => 
                           CARRYB_11_7_port);
   U719 : XNOR2X1 port map( A => n387, B => n501, Y => n934);
   U720 : NAND3X1 port map( A => n859, B => n860, C => n861, Y => n502);
   U721 : XOR2X1 port map( A => CARRYB_12_4_port, B => ab_13_4_port, Y => n811)
                           ;
   U722 : XNOR2X1 port map( A => n504, B => n254, Y => SUMB_14_3_port);
   U723 : INVX1 port map( A => n1051, Y => n505);
   U724 : INVX8 port map( A => B(15), Y => n1051);
   U725 : AND2X2 port map( A => ab_1_11_port, B => ab_0_12_port, Y => n506);
   U726 : INVX1 port map( A => n163, Y => n1040);
   U727 : BUFX4 port map( A => B(9), Y => n507);
   U728 : XOR2X1 port map( A => n94, B => ab_6_4_port, Y => n508);
   U729 : NAND2X1 port map( A => SUMB_5_5_port, B => CARRYB_5_4_port, Y => n509
                           );
   U730 : NAND2X1 port map( A => SUMB_5_5_port, B => ab_6_4_port, Y => n510);
   U731 : NAND2X1 port map( A => CARRYB_5_4_port, B => ab_6_4_port, Y => n511);
   U732 : NAND3X1 port map( A => n511, B => n510, C => n509, Y => 
                           CARRYB_6_4_port);
   U733 : XOR2X1 port map( A => CARRYB_9_9_port, B => ab_10_9_port, Y => n512);
   U734 : XOR2X1 port map( A => SUMB_9_10_port, B => n512, Y => SUMB_10_9_port)
                           ;
   U735 : NAND2X1 port map( A => SUMB_9_10_port, B => CARRYB_9_9_port, Y => 
                           n513);
   U736 : NAND2X1 port map( A => SUMB_9_10_port, B => ab_10_9_port, Y => n514);
   U737 : NAND2X1 port map( A => CARRYB_9_9_port, B => ab_10_9_port, Y => n515)
                           ;
   U738 : NAND3X1 port map( A => n514, B => n513, C => n515, Y => 
                           CARRYB_10_9_port);
   U739 : NAND2X1 port map( A => ab_3_14_port, B => CARRYB_2_14_port, Y => n516
                           );
   U740 : NAND2X1 port map( A => ab_3_14_port, B => ab_2_15_port, Y => n517);
   U741 : NAND2X1 port map( A => CARRYB_2_14_port, B => ab_2_15_port, Y => n518
                           );
   U742 : NAND3X1 port map( A => n516, B => n517, C => n518, Y => 
                           CARRYB_3_14_port);
   U743 : XOR2X1 port map( A => ab_4_14_port, B => ab_3_15_port, Y => n519);
   U744 : XOR2X1 port map( A => n519, B => CARRYB_3_14_port, Y => 
                           SUMB_4_14_port);
   U745 : NAND2X1 port map( A => ab_4_14_port, B => ab_3_15_port, Y => n520);
   U746 : NAND2X1 port map( A => ab_4_14_port, B => CARRYB_3_14_port, Y => n521
                           );
   U747 : NAND2X1 port map( A => ab_3_15_port, B => CARRYB_3_14_port, Y => n522
                           );
   U748 : NAND3X1 port map( A => n520, B => n521, C => n522, Y => 
                           CARRYB_4_14_port);
   U749 : NAND3X1 port map( A => n749, B => n750, C => n751, Y => n523);
   U750 : NAND2X1 port map( A => n527, B => CARRYB_3_1_port, Y => n524);
   U751 : NAND2X1 port map( A => ab_4_1_port, B => n988, Y => n525);
   U752 : NAND2X1 port map( A => n524, B => n525, Y => n616);
   U753 : INVX1 port map( A => ab_4_1_port, Y => n527);
   U754 : INVX8 port map( A => n1012, Y => n1013);
   U755 : INVX4 port map( A => B(13), Y => n1012);
   U756 : BUFX2 port map( A => SUMB_5_4_port, Y => n526);
   U757 : NAND3X1 port map( A => n320, B => n886, C => n887, Y => n528);
   U758 : NAND3X1 port map( A => n950, B => n949, C => n951, Y => n529);
   U759 : XNOR2X1 port map( A => ab_3_2_port, B => n986, Y => n730);
   U760 : INVX2 port map( A => n986, Y => n987);
   U761 : XNOR2X1 port map( A => CARRYB_4_9_port, B => n530, Y => n696);
   U762 : BUFX2 port map( A => A(0), Y => n531);
   U763 : NAND2X1 port map( A => ab_5_3_port, B => n180, Y => n532);
   U764 : NAND2X1 port map( A => ab_5_3_port, B => SUMB_4_4_port, Y => n533);
   U765 : NAND2X1 port map( A => n180, B => SUMB_4_4_port, Y => n534);
   U766 : NAND3X1 port map( A => n532, B => n533, C => n534, Y => 
                           CARRYB_5_3_port);
   U767 : NAND2X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, Y => n535);
   U768 : NAND2X1 port map( A => ab_6_2_port, B => SUMB_5_3_port, Y => n536);
   U769 : NAND2X1 port map( A => CARRYB_5_2_port, B => SUMB_5_3_port, Y => n537
                           );
   U770 : NAND3X1 port map( A => n535, B => n536, C => n537, Y => 
                           CARRYB_6_2_port);
   U771 : AND2X2 port map( A => n1022, B => n1005, Y => n538);
   U772 : INVX1 port map( A => B(8), Y => n1004);
   U773 : INVX4 port map( A => n1004, Y => n1005);
   U774 : XOR2X1 port map( A => CARRYB_4_4_port, B => ab_5_4_port, Y => n539);
   U775 : XOR2X1 port map( A => n469, B => n539, Y => SUMB_5_4_port);
   U776 : NAND2X1 port map( A => SUMB_4_5_port, B => n479, Y => n540);
   U777 : NAND2X1 port map( A => SUMB_4_5_port, B => ab_5_4_port, Y => n541);
   U778 : NAND2X1 port map( A => n479, B => ab_5_4_port, Y => n542);
   U779 : NAND3X1 port map( A => n541, B => n542, C => n540, Y => 
                           CARRYB_5_4_port);
   U780 : XNOR2X1 port map( A => ab_2_3_port, B => n979, Y => n729);
   U781 : NAND3X1 port map( A => n929, B => n928, C => n930, Y => n543);
   U782 : AND2X2 port map( A => n984, B => ab_1_14_port, Y => n961);
   U783 : NAND3X1 port map( A => n879, B => n878, C => n877, Y => n544);
   U784 : NAND2X1 port map( A => SUMB_7_2_port, B => n261, Y => n545);
   U785 : NAND2X1 port map( A => SUMB_7_2_port, B => ab_8_1_port, Y => n546);
   U786 : NAND2X1 port map( A => n261, B => ab_8_1_port, Y => n547);
   U787 : NAND3X1 port map( A => n546, B => n545, C => n547, Y => 
                           CARRYB_8_1_port);
   U788 : BUFX2 port map( A => SUMB_12_1_port, Y => n548);
   U789 : NAND3X1 port map( A => n626, B => n625, C => n627, Y => n549);
   U790 : XOR2X1 port map( A => SUMB_11_1_port, B => ab_12_0_port, Y => n550);
   U791 : XOR2X1 port map( A => n313, B => n550, Y => A1_10_port);
   U792 : NAND2X1 port map( A => CARRYB_11_0_port, B => SUMB_11_1_port, Y => 
                           n551);
   U793 : NAND2X1 port map( A => CARRYB_11_0_port, B => ab_12_0_port, Y => n552
                           );
   U794 : NAND2X1 port map( A => SUMB_11_1_port, B => ab_12_0_port, Y => n553);
   U795 : NAND3X1 port map( A => n553, B => n552, C => n551, Y => 
                           CARRYB_12_0_port);
   U796 : NAND2X1 port map( A => ab_2_7_port, B => n73, Y => n554);
   U797 : NAND2X1 port map( A => SUMB_1_8_port, B => n73, Y => n555);
   U798 : NAND2X1 port map( A => SUMB_1_8_port, B => ab_2_7_port, Y => n556);
   U799 : NAND3X1 port map( A => n556, B => n555, C => n554, Y => 
                           CARRYB_2_7_port);
   U800 : NAND2X1 port map( A => ab_3_6_port, B => n245, Y => n557);
   U801 : NAND2X1 port map( A => SUMB_2_7_port, B => ab_3_6_port, Y => n558);
   U802 : NAND2X1 port map( A => SUMB_2_7_port, B => n245, Y => n559);
   U803 : NAND3X1 port map( A => n557, B => n558, C => n559, Y => 
                           CARRYB_3_6_port);
   U804 : NAND2X1 port map( A => SUMB_1_10_port, B => ab_2_9_port, Y => n560);
   U805 : NAND2X1 port map( A => SUMB_1_10_port, B => n760, Y => n561);
   U806 : NAND2X1 port map( A => n760, B => ab_2_9_port, Y => n562);
   U807 : NAND3X1 port map( A => n561, B => n560, C => n562, Y => 
                           CARRYB_2_9_port);
   U808 : XNOR2X1 port map( A => n569, B => SUMB_9_9_port, Y => SUMB_10_8_port)
                           ;
   U809 : XOR2X1 port map( A => SUMB_7_3_port, B => ab_8_2_port, Y => n563);
   U810 : XOR2X1 port map( A => n322, B => n563, Y => SUMB_8_2_port);
   U811 : NAND2X1 port map( A => SUMB_7_3_port, B => CARRYB_7_2_port, Y => n564
                           );
   U812 : NAND2X1 port map( A => CARRYB_7_2_port, B => ab_8_2_port, Y => n565);
   U813 : NAND2X1 port map( A => SUMB_7_3_port, B => ab_8_2_port, Y => n566);
   U814 : NAND3X1 port map( A => n565, B => n564, C => n566, Y => 
                           CARRYB_8_2_port);
   U815 : XNOR2X1 port map( A => n567, B => n445, Y => SUMB_2_4_port);
   U816 : XNOR2X1 port map( A => n654, B => ab_2_4_port, Y => n567);
   U817 : AND2X2 port map( A => n4, B => n1015, Y => ab_2_14_port);
   U818 : XOR2X1 port map( A => n568, B => n570, Y => n745);
   U819 : XNOR2X1 port map( A => CARRYB_9_8_port, B => ab_10_8_port, Y => n569)
                           ;
   U820 : INVX2 port map( A => CARRYB_11_7_port, Y => n570);
   U821 : NAND2X1 port map( A => SUMB_3_6_port, B => CARRYB_3_5_port, Y => n572
                           );
   U822 : NAND2X1 port map( A => SUMB_3_6_port, B => ab_4_5_port, Y => n573);
   U823 : NAND2X1 port map( A => CARRYB_3_5_port, B => ab_4_5_port, Y => n574);
   U824 : NAND3X1 port map( A => n574, B => n572, C => n573, Y => 
                           CARRYB_4_5_port);
   U825 : XOR2X1 port map( A => n575, B => SUMB_7_8_port, Y => SUMB_8_7_port);
   U826 : NAND2X1 port map( A => ab_7_8_port, B => n466, Y => n576);
   U827 : NAND2X1 port map( A => SUMB_6_9_port, B => ab_7_8_port, Y => n577);
   U828 : NAND2X1 port map( A => n466, B => SUMB_6_9_port, Y => n578);
   U829 : NAND3X1 port map( A => n576, B => n577, C => n578, Y => 
                           CARRYB_7_8_port);
   U830 : NAND2X1 port map( A => ab_8_7_port, B => n394, Y => n579);
   U831 : NAND2X1 port map( A => SUMB_7_8_port, B => ab_8_7_port, Y => n580);
   U832 : NAND2X1 port map( A => SUMB_7_8_port, B => n394, Y => n581);
   U833 : NAND3X1 port map( A => n579, B => n580, C => n581, Y => 
                           CARRYB_8_7_port);
   U834 : NAND3X1 port map( A => n715, B => n717, C => n716, Y => n582);
   U835 : NAND2X1 port map( A => SUMB_6_7_port, B => n300, Y => n583);
   U836 : NAND2X1 port map( A => SUMB_6_7_port, B => ab_7_6_port, Y => n584);
   U837 : NAND2X1 port map( A => n300, B => ab_7_6_port, Y => n585);
   U838 : NAND3X1 port map( A => n585, B => n583, C => n584, Y => 
                           CARRYB_7_6_port);
   U839 : INVX1 port map( A => n1013, Y => n1038);
   U840 : INVX2 port map( A => n981, Y => n982);
   U841 : NOR2X1 port map( A => n1012, B => n655, Y => ab_0_13_port);
   U842 : XOR2X1 port map( A => CARRYB_3_4_port, B => ab_4_4_port, Y => n586);
   U843 : XOR2X1 port map( A => SUMB_3_5_port, B => n586, Y => SUMB_4_4_port);
   U844 : NAND2X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, Y => n587);
   U845 : NAND2X1 port map( A => SUMB_2_6_port, B => ab_3_5_port, Y => n588);
   U846 : NAND2X1 port map( A => CARRYB_2_5_port, B => SUMB_2_6_port, Y => n589
                           );
   U847 : NAND3X1 port map( A => n587, B => n588, C => n589, Y => 
                           CARRYB_3_5_port);
   U848 : NAND2X1 port map( A => ab_4_4_port, B => n549, Y => n590);
   U849 : NAND2X1 port map( A => SUMB_3_5_port, B => ab_4_4_port, Y => n591);
   U850 : NAND2X1 port map( A => SUMB_3_5_port, B => n549, Y => n592);
   U851 : NAND3X1 port map( A => n590, B => n591, C => n592, Y => 
                           CARRYB_4_4_port);
   U852 : INVX1 port map( A => n662, Y => n663);
   U853 : XNOR2X1 port map( A => n803, B => n112, Y => SUMB_5_10_port);
   U854 : XNOR2X1 port map( A => n594, B => SUMB_1_13_port, Y => SUMB_2_12_port
                           );
   U855 : XNOR2X1 port map( A => n802, B => ab_2_12_port, Y => n594);
   U856 : XNOR2X1 port map( A => n595, B => SUMB_14_4_port, Y => SUMB_15_3_port
                           );
   U857 : XOR2X1 port map( A => n219, B => n596, Y => SUMB_3_9_port);
   U858 : NAND2X1 port map( A => SUMB_2_10_port, B => n876, Y => n597);
   U859 : NAND2X1 port map( A => SUMB_2_10_port, B => ab_3_9_port, Y => n598);
   U860 : NAND2X1 port map( A => n876, B => ab_3_9_port, Y => n599);
   U861 : NAND3X1 port map( A => n598, B => n597, C => n599, Y => 
                           CARRYB_3_9_port);
   U862 : NAND3X1 port map( A => n882, B => n881, C => n880, Y => n600);
   U863 : NAND3X1 port map( A => n772, B => n773, C => n774, Y => n601);
   U864 : XOR2X1 port map( A => CARRYB_8_4_port, B => ab_9_4_port, Y => n602);
   U865 : XOR2X1 port map( A => SUMB_8_5_port, B => n602, Y => SUMB_9_4_port);
   U866 : NAND2X1 port map( A => SUMB_8_5_port, B => n544, Y => n603);
   U867 : NAND2X1 port map( A => SUMB_8_5_port, B => ab_9_4_port, Y => n604);
   U868 : NAND2X1 port map( A => n544, B => ab_9_4_port, Y => n605);
   U869 : NAND3X1 port map( A => n605, B => n604, C => n603, Y => 
                           CARRYB_9_4_port);
   U870 : XNOR2X1 port map( A => CARRYB_7_5_port, B => ab_8_5_port, Y => n606);
   U871 : BUFX2 port map( A => SUMB_15_0_port, Y => n607);
   U872 : XOR2X1 port map( A => n86, B => ab_8_0_port, Y => n608);
   U873 : XOR2X1 port map( A => n608, B => n85, Y => A1_6_port);
   U874 : NAND2X1 port map( A => SUMB_7_1_port, B => CARRYB_7_0_port, Y => n609
                           );
   U875 : NAND2X1 port map( A => CARRYB_7_0_port, B => ab_8_0_port, Y => n610);
   U876 : NAND2X1 port map( A => SUMB_7_1_port, B => ab_8_0_port, Y => n611);
   U877 : NAND3X1 port map( A => n611, B => n609, C => n610, Y => 
                           CARRYB_8_0_port);
   U878 : XOR2X1 port map( A => SUMB_6_1_port, B => ab_7_0_port, Y => n612);
   U879 : XOR2X1 port map( A => CARRYB_6_0_port, B => n612, Y => A1_5_port);
   U880 : NAND2X1 port map( A => CARRYB_6_0_port, B => SUMB_6_1_port, Y => n613
                           );
   U881 : NAND2X1 port map( A => CARRYB_6_0_port, B => ab_7_0_port, Y => n614);
   U882 : NAND2X1 port map( A => SUMB_6_1_port, B => ab_7_0_port, Y => n615);
   U883 : NAND3X1 port map( A => n615, B => n613, C => n614, Y => 
                           CARRYB_7_0_port);
   U884 : XOR2X1 port map( A => n616, B => SUMB_3_2_port, Y => SUMB_4_1_port);
   U885 : XOR2X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, Y => n617);
   U886 : XOR2X1 port map( A => n617, B => n360, Y => A1_3_port);
   U887 : NAND2X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, Y => n618);
   U888 : NAND2X1 port map( A => ab_4_1_port, B => SUMB_3_2_port, Y => n619);
   U889 : NAND2X1 port map( A => CARRYB_3_1_port, B => SUMB_3_2_port, Y => n620
                           );
   U890 : NAND3X1 port map( A => n618, B => n619, C => n620, Y => 
                           CARRYB_4_1_port);
   U891 : NAND2X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, Y => n621);
   U892 : NAND2X1 port map( A => ab_5_0_port, B => SUMB_4_1_port, Y => n622);
   U893 : NAND2X1 port map( A => CARRYB_4_0_port, B => SUMB_4_1_port, Y => n623
                           );
   U894 : NAND3X1 port map( A => n621, B => n622, C => n623, Y => 
                           CARRYB_5_0_port);
   U895 : XOR2X1 port map( A => n98, B => n624, Y => SUMB_3_4_port);
   U896 : NAND2X1 port map( A => CARRYB_2_4_port, B => SUMB_2_5_port, Y => n625
                           );
   U897 : NAND2X1 port map( A => SUMB_2_5_port, B => ab_3_4_port, Y => n626);
   U898 : NAND2X1 port map( A => CARRYB_2_4_port, B => ab_3_4_port, Y => n627);
   U899 : NAND3X1 port map( A => n626, B => n625, C => n627, Y => 
                           CARRYB_3_4_port);
   U900 : XOR2X1 port map( A => ab_6_14_port, B => CARRYB_5_14_port, Y => n628)
                           ;
   U901 : XOR2X1 port map( A => n628, B => ab_5_15_port, Y => SUMB_6_14_port);
   U902 : NAND2X1 port map( A => ab_6_14_port, B => CARRYB_5_14_port, Y => n630
                           );
   U903 : NAND2X1 port map( A => ab_6_14_port, B => ab_5_15_port, Y => n631);
   U904 : NAND2X1 port map( A => CARRYB_5_14_port, B => ab_5_15_port, Y => n632
                           );
   U905 : NAND3X1 port map( A => n630, B => n631, C => n632, Y => 
                           CARRYB_6_14_port);
   U906 : NAND2X1 port map( A => ab_7_13_port, B => CARRYB_6_13_port, Y => n633
                           );
   U907 : NAND2X1 port map( A => ab_7_13_port, B => SUMB_6_14_port, Y => n634);
   U908 : NAND2X1 port map( A => CARRYB_6_13_port, B => SUMB_6_14_port, Y => 
                           n635);
   U909 : NAND3X1 port map( A => n633, B => n634, C => n635, Y => 
                           CARRYB_7_13_port);
   U910 : NAND2X1 port map( A => ab_9_11_port, B => CARRYB_8_11_port, Y => n636
                           );
   U911 : NAND2X1 port map( A => SUMB_8_12_port, B => ab_9_11_port, Y => n637);
   U912 : NAND2X1 port map( A => CARRYB_8_11_port, B => SUMB_8_12_port, Y => 
                           n638);
   U913 : NAND3X1 port map( A => n636, B => n637, C => n638, Y => 
                           CARRYB_9_11_port);
   U914 : NAND2X1 port map( A => ab_10_10_port, B => CARRYB_9_10_port, Y => 
                           n639);
   U915 : NAND2X1 port map( A => SUMB_9_11_port, B => ab_10_10_port, Y => n640)
                           ;
   U916 : NAND2X1 port map( A => CARRYB_9_10_port, B => SUMB_9_11_port, Y => 
                           n641);
   U917 : NAND3X1 port map( A => n639, B => n640, C => n641, Y => 
                           CARRYB_10_10_port);
   U918 : XOR2X1 port map( A => n642, B => SUMB_11_9_port, Y => SUMB_12_8_port)
                           ;
   U919 : XOR2X1 port map( A => CARRYB_12_7_port, B => ab_13_7_port, Y => n643)
                           ;
   U920 : NAND2X1 port map( A => ab_12_8_port, B => n20, Y => n644);
   U921 : NAND2X1 port map( A => ab_12_8_port, B => SUMB_11_9_port, Y => n645);
   U922 : NAND2X1 port map( A => n20, B => SUMB_11_9_port, Y => n646);
   U923 : NAND3X1 port map( A => n644, B => n645, C => n646, Y => 
                           CARRYB_12_8_port);
   U924 : NAND2X1 port map( A => ab_13_7_port, B => n523, Y => n647);
   U925 : NAND2X1 port map( A => ab_13_7_port, B => SUMB_12_8_port, Y => n648);
   U926 : NAND2X1 port map( A => n523, B => SUMB_12_8_port, Y => n649);
   U927 : NAND3X1 port map( A => n647, B => n648, C => n649, Y => 
                           CARRYB_13_7_port);
   U928 : XOR2X1 port map( A => CARRYB_7_12_port, B => ab_8_12_port, Y => n650)
                           ;
   U929 : XOR2X1 port map( A => SUMB_7_13_port, B => n650, Y => SUMB_8_12_port)
                           ;
   U930 : NAND2X1 port map( A => SUMB_7_13_port, B => n214, Y => n651);
   U931 : NAND2X1 port map( A => SUMB_7_13_port, B => ab_8_12_port, Y => n652);
   U932 : NAND2X1 port map( A => n214, B => ab_8_12_port, Y => n653);
   U933 : NAND3X1 port map( A => n652, B => n651, C => n653, Y => 
                           CARRYB_8_12_port);
   U934 : AND2X2 port map( A => n962, B => ab_1_4_port, Y => n654);
   U935 : INVX2 port map( A => n907, Y => n984);
   U936 : NAND2X1 port map( A => n49, B => ab_10_3_port, Y => n656);
   U937 : NAND2X1 port map( A => SUMB_9_4_port, B => n49, Y => n657);
   U938 : NAND2X1 port map( A => ab_10_3_port, B => SUMB_9_4_port, Y => n658);
   U939 : NAND3X1 port map( A => n656, B => n657, C => n658, Y => 
                           CARRYB_10_3_port);
   U940 : NAND2X1 port map( A => ab_11_2_port, B => CARRYB_10_2_port, Y => n659
                           );
   U941 : NAND2X1 port map( A => ab_11_2_port, B => SUMB_10_3_port, Y => n660);
   U942 : NAND2X1 port map( A => SUMB_10_3_port, B => CARRYB_10_2_port, Y => 
                           n661);
   U943 : NAND3X1 port map( A => n659, B => n660, C => n661, Y => 
                           CARRYB_11_2_port);
   U944 : INVX2 port map( A => CARRYB_5_5_port, Y => n662);
   U945 : XNOR2X1 port map( A => CARRYB_2_7_port, B => ab_3_7_port, Y => n664);
   U946 : XOR2X1 port map( A => ab_8_10_port, B => CARRYB_7_10_port, Y => n665)
                           ;
   U947 : XOR2X1 port map( A => n665, B => SUMB_7_11_port, Y => SUMB_8_10_port)
                           ;
   U948 : NAND2X1 port map( A => ab_7_11_port, B => CARRYB_6_11_port, Y => n666
                           );
   U949 : NAND2X1 port map( A => ab_7_11_port, B => SUMB_6_12_port, Y => n667);
   U950 : NAND2X1 port map( A => CARRYB_6_11_port, B => SUMB_6_12_port, Y => 
                           n668);
   U951 : NAND3X1 port map( A => n666, B => n667, C => n668, Y => 
                           CARRYB_7_11_port);
   U952 : NAND2X1 port map( A => ab_8_10_port, B => CARRYB_7_10_port, Y => n669
                           );
   U953 : NAND2X1 port map( A => ab_8_10_port, B => SUMB_7_11_port, Y => n670);
   U954 : NAND2X1 port map( A => CARRYB_7_10_port, B => SUMB_7_11_port, Y => 
                           n671);
   U955 : NAND3X1 port map( A => n669, B => n670, C => n671, Y => 
                           CARRYB_8_10_port);
   U956 : XOR2X1 port map( A => ab_9_9_port, B => CARRYB_8_9_port, Y => n672);
   U957 : XOR2X1 port map( A => n672, B => SUMB_8_10_port, Y => SUMB_9_9_port);
   U958 : NAND2X1 port map( A => ab_9_9_port, B => CARRYB_8_9_port, Y => n673);
   U959 : NAND2X1 port map( A => ab_9_9_port, B => SUMB_8_10_port, Y => n674);
   U960 : NAND2X1 port map( A => CARRYB_8_9_port, B => SUMB_8_10_port, Y => 
                           n675);
   U961 : NAND3X1 port map( A => n673, B => n674, C => n675, Y => 
                           CARRYB_9_9_port);
   U962 : NAND2X1 port map( A => ab_10_8_port, B => n55, Y => n676);
   U963 : NAND2X1 port map( A => ab_10_8_port, B => SUMB_9_9_port, Y => n677);
   U964 : NAND2X1 port map( A => n55, B => SUMB_9_9_port, Y => n678);
   U965 : NAND3X1 port map( A => n676, B => n677, C => n678, Y => 
                           CARRYB_10_8_port);
   U966 : NAND2X1 port map( A => ab_14_4_port, B => n268, Y => n679);
   U967 : NAND2X1 port map( A => SUMB_13_5_port, B => ab_14_4_port, Y => n680);
   U968 : NAND2X1 port map( A => SUMB_13_5_port, B => n268, Y => n681);
   U969 : NAND3X1 port map( A => n679, B => n680, C => n681, Y => 
                           CARRYB_14_4_port);
   U970 : NAND2X1 port map( A => ab_15_3_port, B => n392, Y => n682);
   U971 : NAND2X1 port map( A => SUMB_14_4_port, B => ab_15_3_port, Y => n683);
   U972 : NAND2X1 port map( A => SUMB_14_4_port, B => n392, Y => n684);
   U973 : NAND3X1 port map( A => n682, B => n683, C => n684, Y => 
                           CARRYB_15_3_port);
   U974 : XNOR2X1 port map( A => n685, B => SUMB_11_7_port, Y => SUMB_12_6_port
                           );
   U975 : XNOR2X1 port map( A => CARRYB_11_6_port, B => ab_12_6_port, Y => n685
                           );
   U976 : XOR2X1 port map( A => n686, B => n133, Y => SUMB_15_2_port);
   U977 : NAND2X1 port map( A => ab_14_3_port, B => n134, Y => n687);
   U978 : NAND2X1 port map( A => ab_14_3_port, B => SUMB_13_4_port, Y => n688);
   U979 : NAND2X1 port map( A => n134, B => SUMB_13_4_port, Y => n689);
   U980 : NAND3X1 port map( A => n687, B => n688, C => n689, Y => 
                           CARRYB_14_3_port);
   U981 : NAND2X1 port map( A => ab_15_2_port, B => n474, Y => n690);
   U982 : NAND2X1 port map( A => ab_15_2_port, B => SUMB_14_3_port, Y => n691);
   U983 : NAND2X1 port map( A => n474, B => SUMB_14_3_port, Y => n692);
   U984 : NAND3X1 port map( A => n690, B => n692, C => n691, Y => 
                           CARRYB_15_2_port);
   U985 : NAND2X1 port map( A => SUMB_12_5_port, B => n464, Y => n694);
   U986 : NAND2X1 port map( A => n693, B => n811, Y => n695);
   U987 : NAND2X1 port map( A => n695, B => n694, Y => SUMB_13_4_port);
   U988 : INVX1 port map( A => SUMB_12_5_port, Y => n693);
   U989 : XOR2X1 port map( A => n696, B => SUMB_4_10_port, Y => SUMB_5_9_port);
   U990 : NAND2X1 port map( A => ab_5_9_port, B => n502, Y => n697);
   U991 : NAND2X1 port map( A => ab_5_9_port, B => SUMB_4_10_port, Y => n698);
   U992 : NAND2X1 port map( A => SUMB_4_10_port, B => n502, Y => n699);
   U993 : NAND3X1 port map( A => n697, B => n698, C => n699, Y => 
                           CARRYB_5_9_port);
   U994 : NAND2X1 port map( A => SUMB_5_10_port, B => ab_6_9_port, Y => n700);
   U995 : NAND2X1 port map( A => CARRYB_5_9_port, B => ab_6_9_port, Y => n701);
   U996 : NAND2X1 port map( A => SUMB_5_10_port, B => CARRYB_5_9_port, Y => 
                           n702);
   U997 : NAND3X1 port map( A => n700, B => n701, C => n702, Y => 
                           CARRYB_6_9_port);
   U998 : NAND3X1 port map( A => n842, B => n843, C => n844, Y => n703);
   U999 : BUFX2 port map( A => SUMB_13_1_port, Y => n704);
   U1000 : AND2X2 port map( A => SUMB_15_1_port, B => CARRYB_15_0_port, Y => 
                           n955);
   U1001 : INVX2 port map( A => CARRYB_6_2_port, Y => n705);
   U1002 : NAND2X1 port map( A => ab_11_6_port, B => n88, Y => n706);
   U1003 : NAND2X1 port map( A => SUMB_10_7_port, B => ab_11_6_port, Y => n707)
                           ;
   U1004 : NAND2X1 port map( A => SUMB_10_7_port, B => n88, Y => n708);
   U1005 : NAND3X1 port map( A => n706, B => n707, C => n708, Y => 
                           CARRYB_11_6_port);
   U1006 : NAND2X1 port map( A => ab_12_5_port, B => n154, Y => n709);
   U1007 : NAND2X1 port map( A => SUMB_11_6_port, B => ab_12_5_port, Y => n710)
                           ;
   U1008 : NAND2X1 port map( A => n154, B => SUMB_11_6_port, Y => n711);
   U1009 : NAND3X1 port map( A => n709, B => n710, C => n711, Y => 
                           CARRYB_12_5_port);
   U1010 : NAND2X1 port map( A => n160, B => n183, Y => n712);
   U1011 : NAND2X1 port map( A => SUMB_1_13_port, B => n183, Y => n713);
   U1012 : NAND2X1 port map( A => SUMB_1_13_port, B => n160, Y => n714);
   U1013 : NAND3X1 port map( A => n712, B => n713, C => n714, Y => 
                           CARRYB_2_12_port);
   U1014 : NAND2X1 port map( A => ab_3_11_port, B => CARRYB_2_11_port, Y => 
                           n715);
   U1015 : NAND2X1 port map( A => SUMB_2_12_port, B => ab_3_11_port, Y => n716)
                           ;
   U1016 : NAND2X1 port map( A => SUMB_2_12_port, B => CARRYB_2_11_port, Y => 
                           n717);
   U1017 : NAND3X1 port map( A => n715, B => n716, C => n717, Y => 
                           CARRYB_3_11_port);
   U1018 : XNOR2X1 port map( A => n718, B => SUMB_9_8_port, Y => SUMB_10_7_port
                           );
   U1019 : XNOR2X1 port map( A => ab_10_7_port, B => CARRYB_9_7_port, Y => n718
                           );
   U1020 : NAND2X1 port map( A => n7, B => SUMB_9_2_port, Y => n719);
   U1021 : NAND2X1 port map( A => CARRYB_9_1_port, B => ab_10_1_port, Y => n720
                           );
   U1022 : NAND2X1 port map( A => SUMB_9_2_port, B => ab_10_1_port, Y => n721);
   U1023 : NAND3X1 port map( A => n720, B => n721, C => n719, Y => 
                           CARRYB_10_1_port);
   U1024 : NAND2X1 port map( A => SUMB_6_2_port, B => CARRYB_6_1_port, Y => 
                           n722);
   U1025 : NAND2X1 port map( A => CARRYB_6_1_port, B => ab_7_1_port, Y => n723)
                           ;
   U1026 : NAND2X1 port map( A => SUMB_6_2_port, B => ab_7_1_port, Y => n724);
   U1027 : NAND3X1 port map( A => n724, B => n722, C => n723, Y => 
                           CARRYB_7_1_port);
   U1028 : XOR2X1 port map( A => CARRYB_4_1_port, B => ab_5_1_port, Y => n725);
   U1029 : XOR2X1 port map( A => SUMB_4_2_port, B => n725, Y => SUMB_5_1_port);
   U1030 : NAND2X1 port map( A => SUMB_4_2_port, B => CARRYB_4_1_port, Y => 
                           n726);
   U1031 : NAND2X1 port map( A => SUMB_4_2_port, B => ab_5_1_port, Y => n727);
   U1032 : NAND2X1 port map( A => CARRYB_4_1_port, B => ab_5_1_port, Y => n728)
                           ;
   U1033 : NAND3X1 port map( A => n727, B => n728, C => n726, Y => 
                           CARRYB_5_1_port);
   U1034 : XOR2X1 port map( A => n729, B => SUMB_1_4_port, Y => SUMB_2_3_port);
   U1035 : XOR2X1 port map( A => n730, B => SUMB_2_3_port, Y => SUMB_3_2_port);
   U1036 : NAND2X1 port map( A => ab_2_3_port, B => n959, Y => n731);
   U1037 : NAND2X1 port map( A => ab_2_3_port, B => SUMB_1_4_port, Y => n732);
   U1038 : NAND2X1 port map( A => n959, B => SUMB_1_4_port, Y => n733);
   U1039 : NAND3X1 port map( A => n731, B => n732, C => n733, Y => 
                           CARRYB_2_3_port);
   U1040 : NAND2X1 port map( A => ab_3_2_port, B => n987, Y => n734);
   U1041 : NAND2X1 port map( A => ab_3_2_port, B => SUMB_2_3_port, Y => n735);
   U1042 : NAND2X1 port map( A => n987, B => SUMB_2_3_port, Y => n736);
   U1043 : NAND3X1 port map( A => n734, B => n735, C => n736, Y => 
                           CARRYB_3_2_port);
   U1044 : XNOR2X1 port map( A => CARRYB_3_7_port, B => ab_4_7_port, Y => n737)
                           ;
   U1045 : NAND2X1 port map( A => SUMB_6_4_port, B => n529, Y => n738);
   U1046 : NAND2X1 port map( A => SUMB_6_4_port, B => ab_7_3_port, Y => n739);
   U1047 : NAND2X1 port map( A => n529, B => ab_7_3_port, Y => n740);
   U1048 : NAND3X1 port map( A => n739, B => n740, C => n738, Y => 
                           CARRYB_7_3_port);
   U1049 : XOR2X1 port map( A => n528, B => ab_13_1_port, Y => n837);
   U1050 : XOR2X1 port map( A => SUMB_14_5_port, B => n741, Y => SUMB_15_4_port
                           );
   U1051 : NAND2X1 port map( A => SUMB_14_5_port, B => n270, Y => n742);
   U1052 : NAND2X1 port map( A => SUMB_14_5_port, B => ab_15_4_port, Y => n743)
                           ;
   U1053 : NAND2X1 port map( A => n270, B => ab_15_4_port, Y => n744);
   U1054 : NAND3X1 port map( A => n744, B => n742, C => n743, Y => 
                           CARRYB_15_4_port);
   U1055 : XOR2X1 port map( A => n745, B => SUMB_11_8_port, Y => SUMB_12_7_port
                           );
   U1056 : NAND2X1 port map( A => ab_11_8_port, B => CARRYB_10_8_port, Y => 
                           n746);
   U1057 : NAND2X1 port map( A => ab_11_8_port, B => SUMB_10_9_port, Y => n747)
                           ;
   U1058 : NAND2X1 port map( A => CARRYB_10_8_port, B => SUMB_10_9_port, Y => 
                           n748);
   U1059 : NAND3X1 port map( A => n746, B => n747, C => n748, Y => 
                           CARRYB_11_8_port);
   U1060 : NAND2X1 port map( A => ab_12_7_port, B => n571, Y => n749);
   U1061 : NAND2X1 port map( A => SUMB_11_8_port, B => ab_12_7_port, Y => n750)
                           ;
   U1062 : NAND2X1 port map( A => n571, B => SUMB_11_8_port, Y => n751);
   U1063 : NAND3X1 port map( A => n749, B => n750, C => n751, Y => 
                           CARRYB_12_7_port);
   U1064 : XOR2X1 port map( A => ab_7_12_port, B => n239, Y => n752);
   U1065 : XOR2X1 port map( A => n752, B => SUMB_6_13_port, Y => SUMB_7_12_port
                           );
   U1066 : XOR2X1 port map( A => CARRYB_7_11_port, B => ab_8_11_port, Y => n753
                           );
   U1067 : XOR2X1 port map( A => n753, B => SUMB_7_12_port, Y => SUMB_8_11_port
                           );
   U1068 : NAND2X1 port map( A => ab_7_12_port, B => n239, Y => n754);
   U1069 : NAND2X1 port map( A => ab_7_12_port, B => SUMB_6_13_port, Y => n755)
                           ;
   U1070 : NAND2X1 port map( A => n239, B => SUMB_6_13_port, Y => n756);
   U1071 : NAND3X1 port map( A => n754, B => n755, C => n756, Y => 
                           CARRYB_7_12_port);
   U1072 : NAND2X1 port map( A => ab_8_11_port, B => CARRYB_7_11_port, Y => 
                           n757);
   U1073 : NAND2X1 port map( A => ab_8_11_port, B => SUMB_7_12_port, Y => n758)
                           ;
   U1074 : NAND2X1 port map( A => CARRYB_7_11_port, B => SUMB_7_12_port, Y => 
                           n759);
   U1075 : NAND3X1 port map( A => n757, B => n758, C => n759, Y => 
                           CARRYB_8_11_port);
   U1076 : AND2X2 port map( A => ab_0_10_port, B => ab_1_9_port, Y => n760);
   U1077 : XOR2X1 port map( A => A(15), B => n505, Y => n761);
   U1078 : XOR2X1 port map( A => n607, B => n761, Y => A1_13_port);
   U1079 : NAND2X1 port map( A => SUMB_15_0_port, B => A(15), Y => n762);
   U1080 : NAND2X1 port map( A => SUMB_15_0_port, B => n505, Y => n763);
   U1081 : NAND2X1 port map( A => A(15), B => n505, Y => n764);
   U1082 : NAND3X1 port map( A => n764, B => n763, C => n762, Y => A2_14_port);
   U1083 : NAND2X1 port map( A => ab_11_3_port, B => n159, Y => n765);
   U1084 : NAND2X1 port map( A => SUMB_10_4_port, B => ab_11_3_port, Y => n766)
                           ;
   U1085 : NAND2X1 port map( A => n159, B => SUMB_10_4_port, Y => n767);
   U1086 : NAND3X1 port map( A => n765, B => n766, C => n767, Y => 
                           CARRYB_11_3_port);
   U1087 : NAND2X1 port map( A => n95, B => ab_12_2_port, Y => n768);
   U1088 : NAND2X1 port map( A => SUMB_11_3_port, B => n95, Y => n769);
   U1089 : NAND2X1 port map( A => SUMB_11_3_port, B => ab_12_2_port, Y => n770)
                           ;
   U1090 : NAND3X1 port map( A => n768, B => n770, C => n769, Y => 
                           CARRYB_12_2_port);
   U1091 : XOR2X1 port map( A => SUMB_4_8_port, B => n771, Y => SUMB_5_7_port);
   U1092 : NAND2X1 port map( A => ab_4_8_port, B => n390, Y => n772);
   U1093 : NAND2X1 port map( A => SUMB_3_9_port, B => ab_4_8_port, Y => n773);
   U1094 : NAND2X1 port map( A => n390, B => SUMB_3_9_port, Y => n774);
   U1095 : NAND3X1 port map( A => n772, B => n773, C => n774, Y => 
                           CARRYB_4_8_port);
   U1096 : NAND2X1 port map( A => ab_5_7_port, B => n377, Y => n775);
   U1097 : NAND2X1 port map( A => SUMB_4_8_port, B => ab_5_7_port, Y => n776);
   U1098 : NAND2X1 port map( A => SUMB_4_8_port, B => n377, Y => n777);
   U1099 : NAND3X1 port map( A => n775, B => n776, C => n777, Y => 
                           CARRYB_5_7_port);
   U1100 : INVX1 port map( A => n1007, Y => n1041);
   U1101 : NAND2X1 port map( A => ab_9_7_port, B => n467, Y => n778);
   U1102 : NAND2X1 port map( A => SUMB_8_8_port, B => ab_9_7_port, Y => n779);
   U1103 : NAND2X1 port map( A => n467, B => SUMB_8_8_port, Y => n780);
   U1104 : NAND3X1 port map( A => n778, B => n779, C => n780, Y => 
                           CARRYB_9_7_port);
   U1105 : NAND2X1 port map( A => n391, B => ab_10_6_port, Y => n781);
   U1106 : NAND2X1 port map( A => SUMB_9_7_port, B => n391, Y => n782);
   U1107 : NAND2X1 port map( A => SUMB_9_7_port, B => ab_10_6_port, Y => n783);
   U1108 : NAND3X1 port map( A => n781, B => n782, C => n783, Y => 
                           CARRYB_10_6_port);
   U1109 : INVX1 port map( A => n1011, Y => n1039);
   U1110 : NAND2X1 port map( A => ab_3_7_port, B => n396, Y => n784);
   U1111 : NAND2X1 port map( A => SUMB_2_8_port, B => ab_3_7_port, Y => n785);
   U1112 : NAND2X1 port map( A => SUMB_2_8_port, B => n396, Y => n786);
   U1113 : NAND3X1 port map( A => n784, B => n785, C => n786, Y => 
                           CARRYB_3_7_port);
   U1114 : NAND2X1 port map( A => n446, B => ab_4_6_port, Y => n787);
   U1115 : NAND2X1 port map( A => SUMB_3_7_port, B => ab_4_6_port, Y => n788);
   U1116 : NAND2X1 port map( A => SUMB_3_7_port, B => n446, Y => n789);
   U1117 : NAND3X1 port map( A => n787, B => n789, C => n788, Y => 
                           CARRYB_4_6_port);
   U1118 : NAND2X1 port map( A => SUMB_1_9_port, B => n415, Y => n790);
   U1119 : NAND2X1 port map( A => ab_2_8_port, B => n415, Y => n791);
   U1120 : NAND2X1 port map( A => SUMB_1_9_port, B => ab_2_8_port, Y => n792);
   U1121 : NAND2X1 port map( A => ab_10_5_port, B => n93, Y => n793);
   U1122 : NAND2X1 port map( A => SUMB_9_6_port, B => ab_10_5_port, Y => n794);
   U1123 : NAND2X1 port map( A => SUMB_9_6_port, B => n93, Y => n795);
   U1124 : NAND3X1 port map( A => n794, B => n793, C => n795, Y => 
                           CARRYB_10_5_port);
   U1125 : NAND2X1 port map( A => ab_11_4_port, B => n971, Y => n796);
   U1126 : NAND2X1 port map( A => SUMB_10_5_port, B => ab_11_4_port, Y => n797)
                           ;
   U1127 : NAND2X1 port map( A => SUMB_10_5_port, B => n971, Y => n798);
   U1128 : NAND3X1 port map( A => n796, B => n797, C => n798, Y => 
                           CARRYB_11_4_port);
   U1129 : NAND2X1 port map( A => SUMB_8_7_port, B => CARRYB_8_6_port, Y => 
                           n799);
   U1130 : NAND2X1 port map( A => SUMB_8_7_port, B => ab_9_6_port, Y => n800);
   U1131 : NAND2X1 port map( A => n45, B => ab_9_6_port, Y => n801);
   U1132 : NAND3X1 port map( A => n801, B => n799, C => n800, Y => 
                           CARRYB_9_6_port);
   U1133 : AND2X2 port map( A => ab_0_13_port, B => ab_1_12_port, Y => n802);
   U1134 : XOR2X1 port map( A => n981, B => n804, Y => n883);
   U1135 : NAND2X1 port map( A => ab_9_8_port, B => n236, Y => n805);
   U1136 : NAND2X1 port map( A => SUMB_8_9_port, B => ab_9_8_port, Y => n806);
   U1137 : NAND2X1 port map( A => n236, B => SUMB_8_9_port, Y => n807);
   U1138 : NAND3X1 port map( A => n805, B => n806, C => n807, Y => 
                           CARRYB_9_8_port);
   U1139 : NAND2X1 port map( A => ab_10_7_port, B => n272, Y => n808);
   U1140 : NAND2X1 port map( A => SUMB_9_8_port, B => ab_10_7_port, Y => n809);
   U1141 : NAND2X1 port map( A => SUMB_9_8_port, B => n272, Y => n810);
   U1142 : NAND3X1 port map( A => n808, B => n809, C => n810, Y => 
                           CARRYB_10_7_port);
   U1143 : NAND2X1 port map( A => SUMB_12_5_port, B => n703, Y => n812);
   U1144 : NAND2X1 port map( A => SUMB_12_5_port, B => ab_13_4_port, Y => n813)
                           ;
   U1145 : NAND2X1 port map( A => n703, B => ab_13_4_port, Y => n814);
   U1146 : NAND3X1 port map( A => n813, B => n812, C => n814, Y => 
                           CARRYB_13_4_port);
   U1147 : NAND2X1 port map( A => SUMB_7_9_port, B => n480, Y => n815);
   U1148 : NAND2X1 port map( A => SUMB_7_9_port, B => ab_8_8_port, Y => n816);
   U1149 : NAND2X1 port map( A => n480, B => ab_8_8_port, Y => n817);
   U1150 : NAND3X1 port map( A => n816, B => n815, C => n817, Y => 
                           CARRYB_8_8_port);
   U1151 : NAND2X1 port map( A => ab_4_10_port, B => CARRYB_3_10_port, Y => 
                           n818);
   U1152 : NAND2X1 port map( A => ab_4_10_port, B => SUMB_3_11_port, Y => n819)
                           ;
   U1153 : NAND2X1 port map( A => CARRYB_3_10_port, B => SUMB_3_11_port, Y => 
                           n820);
   U1154 : NAND2X1 port map( A => n77, B => ab_5_10_port, Y => n821);
   U1155 : NAND2X1 port map( A => ab_5_10_port, B => n112, Y => n822);
   U1156 : NAND2X1 port map( A => n77, B => n112, Y => n823);
   U1157 : NAND3X1 port map( A => n821, B => n822, C => n823, Y => 
                           CARRYB_5_10_port);
   U1158 : NAND2X1 port map( A => ab_12_6_port, B => n273, Y => n824);
   U1159 : NAND2X1 port map( A => SUMB_11_7_port, B => ab_12_6_port, Y => n825)
                           ;
   U1160 : NAND2X1 port map( A => SUMB_11_7_port, B => n273, Y => n826);
   U1161 : NAND3X1 port map( A => n824, B => n825, C => n826, Y => 
                           CARRYB_12_6_port);
   U1162 : NAND2X1 port map( A => ab_13_5_port, B => n82, Y => n827);
   U1163 : NAND2X1 port map( A => SUMB_12_6_port, B => ab_13_5_port, Y => n828)
                           ;
   U1164 : NAND2X1 port map( A => SUMB_12_6_port, B => n82, Y => n829);
   U1165 : XOR2X1 port map( A => n345, B => ab_6_11_port, Y => n830);
   U1166 : XOR2X1 port map( A => n830, B => SUMB_5_12_port, Y => SUMB_6_11_port
                           );
   U1167 : NAND2X1 port map( A => SUMB_5_12_port, B => n345, Y => n831);
   U1168 : NAND2X1 port map( A => SUMB_5_12_port, B => ab_6_11_port, Y => n832)
                           ;
   U1169 : NAND2X1 port map( A => n345, B => ab_6_11_port, Y => n833);
   U1170 : NAND3X1 port map( A => n832, B => n831, C => n833, Y => 
                           CARRYB_6_11_port);
   U1171 : NAND2X1 port map( A => SUMB_7_10_port, B => CARRYB_7_9_port, Y => 
                           n834);
   U1172 : NAND2X1 port map( A => CARRYB_7_9_port, B => ab_8_9_port, Y => n835)
                           ;
   U1173 : NAND2X1 port map( A => SUMB_7_10_port, B => ab_8_9_port, Y => n836);
   U1174 : NAND3X1 port map( A => n835, B => n834, C => n836, Y => 
                           CARRYB_8_9_port);
   U1175 : INVX1 port map( A => n1015, Y => n1037);
   U1176 : NAND2X1 port map( A => CARRYB_12_1_port, B => SUMB_12_2_port, Y => 
                           n838);
   U1177 : NAND2X1 port map( A => SUMB_12_2_port, B => ab_13_1_port, Y => n839)
                           ;
   U1178 : NAND2X1 port map( A => CARRYB_12_1_port, B => ab_13_1_port, Y => 
                           n840);
   U1179 : NAND3X1 port map( A => n839, B => n838, C => n840, Y => 
                           CARRYB_13_1_port);
   U1180 : INVX2 port map( A => CARRYB_3_6_port, Y => n841);
   U1181 : NAND2X1 port map( A => ab_12_4_port, B => n369, Y => n842);
   U1182 : NAND2X1 port map( A => SUMB_11_5_port, B => ab_12_4_port, Y => n843)
                           ;
   U1183 : NAND2X1 port map( A => SUMB_11_5_port, B => n369, Y => n844);
   U1184 : NAND3X1 port map( A => n842, B => n843, C => n844, Y => 
                           CARRYB_12_4_port);
   U1185 : NAND2X1 port map( A => CARRYB_12_3_port, B => ab_13_3_port, Y => 
                           n845);
   U1186 : NAND2X1 port map( A => ab_13_3_port, B => SUMB_12_4_port, Y => n846)
                           ;
   U1187 : NAND2X1 port map( A => SUMB_12_4_port, B => CARRYB_12_3_port, Y => 
                           n847);
   U1188 : NAND2X1 port map( A => SUMB_3_13_port, B => n346, Y => n848);
   U1189 : NAND2X1 port map( A => SUMB_3_13_port, B => ab_4_12_port, Y => n849)
                           ;
   U1190 : NAND2X1 port map( A => n346, B => ab_4_12_port, Y => n850);
   U1191 : NAND3X1 port map( A => n849, B => n848, C => n850, Y => 
                           CARRYB_4_12_port);
   U1192 : XOR2X1 port map( A => ab_5_11_port, B => CARRYB_4_11_port, Y => n851
                           );
   U1193 : XOR2X1 port map( A => n851, B => SUMB_4_12_port, Y => SUMB_5_11_port
                           );
   U1194 : XOR2X1 port map( A => n852, B => n18, Y => SUMB_6_10_port);
   U1195 : NAND2X1 port map( A => ab_5_11_port, B => n249, Y => n853);
   U1196 : NAND2X1 port map( A => SUMB_4_12_port, B => ab_5_11_port, Y => n854)
                           ;
   U1197 : NAND2X1 port map( A => SUMB_4_12_port, B => n249, Y => n855);
   U1198 : NAND2X1 port map( A => ab_6_10_port, B => CARRYB_5_10_port, Y => 
                           n856);
   U1199 : NAND2X1 port map( A => ab_6_10_port, B => SUMB_5_11_port, Y => n857)
                           ;
   U1200 : NAND2X1 port map( A => CARRYB_5_10_port, B => SUMB_5_11_port, Y => 
                           n858);
   U1201 : NAND3X1 port map( A => n856, B => n857, C => n858, Y => 
                           CARRYB_6_10_port);
   U1202 : NAND2X1 port map( A => ab_4_9_port, B => CARRYB_3_9_port, Y => n859)
                           ;
   U1203 : NAND2X1 port map( A => SUMB_3_10_port, B => ab_4_9_port, Y => n860);
   U1204 : NAND2X1 port map( A => CARRYB_3_9_port, B => SUMB_3_10_port, Y => 
                           n861);
   U1205 : NAND3X1 port map( A => n860, B => n859, C => n861, Y => 
                           CARRYB_4_9_port);
   U1206 : NAND2X1 port map( A => ab_5_8_port, B => n601, Y => n862);
   U1207 : NAND2X1 port map( A => SUMB_4_9_port, B => ab_5_8_port, Y => n863);
   U1208 : NAND2X1 port map( A => SUMB_4_9_port, B => n601, Y => n864);
   U1209 : NAND3X1 port map( A => n862, B => n863, C => n864, Y => 
                           CARRYB_5_8_port);
   U1210 : NAND2X1 port map( A => ab_8_6_port, B => n318, Y => n865);
   U1211 : NAND2X1 port map( A => SUMB_7_7_port, B => ab_8_6_port, Y => n866);
   U1212 : NAND2X1 port map( A => SUMB_7_7_port, B => n318, Y => n867);
   U1213 : NAND3X1 port map( A => n865, B => n866, C => n867, Y => 
                           CARRYB_8_6_port);
   U1214 : NAND2X1 port map( A => ab_9_5_port, B => n600, Y => n868);
   U1215 : NAND2X1 port map( A => ab_9_5_port, B => SUMB_8_6_port, Y => n869);
   U1216 : NAND2X1 port map( A => n600, B => SUMB_8_6_port, Y => n870);
   U1217 : NAND3X1 port map( A => n868, B => n869, C => n870, Y => 
                           CARRYB_9_5_port);
   U1218 : XOR2X1 port map( A => n386, B => ab_14_0_port, Y => n871);
   U1219 : XOR2X1 port map( A => n704, B => n871, Y => A1_12_port);
   U1220 : NAND2X1 port map( A => SUMB_13_1_port, B => CARRYB_13_0_port, Y => 
                           n872);
   U1221 : NAND2X1 port map( A => SUMB_13_1_port, B => ab_14_0_port, Y => n873)
                           ;
   U1222 : NAND2X1 port map( A => CARRYB_13_0_port, B => ab_14_0_port, Y => 
                           n874);
   U1223 : NAND3X1 port map( A => n874, B => n872, C => n873, Y => 
                           CARRYB_14_0_port);
   U1224 : NAND2X1 port map( A => SUMB_7_5_port, B => n543, Y => n877);
   U1225 : NAND2X1 port map( A => SUMB_7_5_port, B => ab_8_4_port, Y => n878);
   U1226 : NAND2X1 port map( A => n543, B => ab_8_4_port, Y => n879);
   U1227 : NAND3X1 port map( A => n879, B => n877, C => n878, Y => 
                           CARRYB_8_4_port);
   U1228 : NAND2X1 port map( A => SUMB_7_6_port, B => n278, Y => n880);
   U1229 : NAND2X1 port map( A => SUMB_7_6_port, B => ab_8_5_port, Y => n881);
   U1230 : NAND2X1 port map( A => n278, B => ab_8_5_port, Y => n882);
   U1231 : NAND3X1 port map( A => n882, B => n881, C => n880, Y => 
                           CARRYB_8_5_port);
   U1232 : XOR2X1 port map( A => ab_13_0_port, B => n388, Y => n884);
   U1233 : XOR2X1 port map( A => n884, B => n548, Y => A1_11_port);
   U1234 : NAND2X1 port map( A => ab_12_1_port, B => n982, Y => n885);
   U1235 : NAND2X1 port map( A => SUMB_11_2_port, B => ab_12_1_port, Y => n886)
                           ;
   U1236 : NAND2X1 port map( A => n982, B => SUMB_11_2_port, Y => n887);
   U1237 : NAND3X1 port map( A => n885, B => n887, C => n886, Y => 
                           CARRYB_12_1_port);
   U1238 : NAND2X1 port map( A => CARRYB_12_0_port, B => ab_13_0_port, Y => 
                           n888);
   U1239 : NAND2X1 port map( A => ab_13_0_port, B => SUMB_12_1_port, Y => n889)
                           ;
   U1240 : NAND2X1 port map( A => CARRYB_12_0_port, B => SUMB_12_1_port, Y => 
                           n890);
   U1241 : NAND3X1 port map( A => n889, B => n890, C => n888, Y => 
                           CARRYB_13_0_port);
   U1242 : NAND2X1 port map( A => n538, B => n301, Y => n891);
   U1243 : NAND2X1 port map( A => SUMB_2_9_port, B => n538, Y => n892);
   U1244 : NAND2X1 port map( A => SUMB_2_9_port, B => n301, Y => n893);
   U1245 : NAND3X1 port map( A => n891, B => n892, C => n893, Y => 
                           CARRYB_3_8_port);
   U1246 : NAND2X1 port map( A => n475, B => ab_4_7_port, Y => n894);
   U1247 : NAND2X1 port map( A => ab_4_7_port, B => SUMB_3_8_port, Y => n895);
   U1248 : NAND2X1 port map( A => SUMB_3_8_port, B => n475, Y => n896);
   U1249 : NAND3X1 port map( A => n894, B => n896, C => n895, Y => 
                           CARRYB_4_7_port);
   U1250 : XOR2X1 port map( A => SUMB_6_8_port, B => n897, Y => SUMB_7_7_port);
   U1251 : NAND2X1 port map( A => ab_6_8_port, B => n393, Y => n898);
   U1252 : NAND2X1 port map( A => SUMB_5_9_port, B => ab_6_8_port, Y => n899);
   U1253 : NAND2X1 port map( A => SUMB_5_9_port, B => n393, Y => n900);
   U1254 : NAND3X1 port map( A => n898, B => n899, C => n900, Y => 
                           CARRYB_6_8_port);
   U1255 : NAND2X1 port map( A => n44, B => ab_7_7_port, Y => n901);
   U1256 : NAND2X1 port map( A => SUMB_6_8_port, B => ab_7_7_port, Y => n902);
   U1257 : NAND2X1 port map( A => SUMB_6_8_port, B => n256, Y => n903);
   U1258 : NAND3X1 port map( A => n901, B => n902, C => n903, Y => 
                           CARRYB_7_7_port);
   U1259 : INVX1 port map( A => n507, Y => n1042);
   U1260 : AND2X2 port map( A => ab_1_6_port, B => ab_0_7_port, Y => n904);
   U1261 : INVX2 port map( A => n1002, Y => n1003);
   U1262 : INVX2 port map( A => B(7), Y => n1002);
   U1263 : INVX1 port map( A => n905, Y => n1043);
   U1264 : INVX4 port map( A => n1000, Y => n969);
   U1265 : AND2X2 port map( A => ab_1_7_port, B => ab_0_8_port, Y => n906);
   U1266 : NAND2X1 port map( A => n655, B => B(15), Y => n907);
   U1267 : NAND2X1 port map( A => ab_3_12_port, B => n271, Y => n908);
   U1268 : NAND2X1 port map( A => SUMB_2_13_port, B => ab_3_12_port, Y => n909)
                           ;
   U1269 : NAND2X1 port map( A => n271, B => SUMB_2_13_port, Y => n910);
   U1270 : NAND3X1 port map( A => n908, B => n909, C => n910, Y => 
                           CARRYB_3_12_port);
   U1271 : NAND2X1 port map( A => ab_4_11_port, B => n582, Y => n911);
   U1272 : NAND2X1 port map( A => SUMB_3_12_port, B => ab_4_11_port, Y => n912)
                           ;
   U1273 : NAND2X1 port map( A => SUMB_3_12_port, B => n582, Y => n913);
   U1274 : NAND3X1 port map( A => n911, B => n912, C => n913, Y => 
                           CARRYB_4_11_port);
   U1275 : XOR2X1 port map( A => SUMB_1_14_port, B => n914, Y => SUMB_2_13_port
                           );
   U1276 : NAND2X1 port map( A => SUMB_1_14_port, B => ab_2_13_port, Y => n915)
                           ;
   U1277 : NAND2X1 port map( A => SUMB_1_14_port, B => n246, Y => n916);
   U1278 : NAND2X1 port map( A => ab_2_13_port, B => n246, Y => n917);
   U1279 : NAND3X1 port map( A => n916, B => n915, C => n917, Y => 
                           CARRYB_2_13_port);
   U1280 : XOR2X1 port map( A => n918, B => n76, Y => SUMB_14_1_port);
   U1281 : NAND2X1 port map( A => ab_13_2_port, B => n398, Y => n919);
   U1282 : NAND2X1 port map( A => SUMB_12_3_port, B => ab_13_2_port, Y => n920)
                           ;
   U1283 : NAND2X1 port map( A => SUMB_12_3_port, B => n398, Y => n921);
   U1284 : NAND3X1 port map( A => n919, B => n921, C => n920, Y => 
                           CARRYB_13_2_port);
   U1285 : NAND2X1 port map( A => ab_14_1_port, B => n87, Y => n922);
   U1286 : NAND2X1 port map( A => SUMB_13_2_port, B => ab_14_1_port, Y => n923)
                           ;
   U1287 : NAND2X1 port map( A => SUMB_13_2_port, B => n87, Y => n924);
   U1288 : NAND3X1 port map( A => n922, B => n923, C => n924, Y => 
                           CARRYB_14_1_port);
   U1289 : NAND2X1 port map( A => ab_6_5_port, B => n663, Y => n925);
   U1290 : NAND2X1 port map( A => SUMB_5_6_port, B => ab_6_5_port, Y => n926);
   U1291 : NAND2X1 port map( A => SUMB_5_6_port, B => n663, Y => n927);
   U1292 : NAND3X1 port map( A => n926, B => n925, C => n927, Y => 
                           CARRYB_6_5_port);
   U1293 : NAND2X1 port map( A => n14, B => ab_7_4_port, Y => n928);
   U1294 : NAND2X1 port map( A => SUMB_6_5_port, B => ab_7_4_port, Y => n929);
   U1295 : NAND2X1 port map( A => n14, B => SUMB_6_5_port, Y => n930);
   U1296 : NAND3X1 port map( A => n928, B => n929, C => n930, Y => 
                           CARRYB_7_4_port);
   U1297 : NAND2X1 port map( A => SUMB_9_3_port, B => n15, Y => n931);
   U1298 : NAND2X1 port map( A => SUMB_9_3_port, B => ab_10_2_port, Y => n932);
   U1299 : NAND2X1 port map( A => n15, B => ab_10_2_port, Y => n933);
   U1300 : NAND3X1 port map( A => n932, B => n931, C => n933, Y => 
                           CARRYB_10_2_port);
   U1301 : XOR2X1 port map( A => ab_5_2_port, B => n164, Y => n935);
   U1302 : XOR2X1 port map( A => n935, B => n321, Y => SUMB_5_2_port);
   U1303 : NAND2X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, Y => n936)
                           ;
   U1304 : NAND2X1 port map( A => ab_4_3_port, B => SUMB_3_4_port, Y => n937);
   U1305 : NAND2X1 port map( A => CARRYB_3_3_port, B => SUMB_3_4_port, Y => 
                           n938);
   U1306 : NAND3X1 port map( A => n936, B => n937, C => n938, Y => 
                           CARRYB_4_3_port);
   U1307 : NAND2X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, Y => n939)
                           ;
   U1308 : NAND2X1 port map( A => ab_5_2_port, B => SUMB_4_3_port, Y => n940);
   U1309 : NAND2X1 port map( A => CARRYB_4_2_port, B => SUMB_4_3_port, Y => 
                           n941);
   U1310 : NAND3X1 port map( A => n939, B => n940, C => n941, Y => 
                           CARRYB_5_2_port);
   U1311 : NAND2X1 port map( A => ab_2_4_port, B => n654, Y => n942);
   U1312 : NAND2X1 port map( A => ab_2_4_port, B => SUMB_1_5_port, Y => n943);
   U1313 : NAND2X1 port map( A => n654, B => SUMB_1_5_port, Y => n944);
   U1314 : NAND3X1 port map( A => n942, B => n943, C => n944, Y => 
                           CARRYB_2_4_port);
   U1315 : NAND2X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, Y => n945)
                           ;
   U1316 : NAND2X1 port map( A => ab_3_3_port, B => SUMB_2_4_port, Y => n946);
   U1317 : NAND2X1 port map( A => CARRYB_2_3_port, B => SUMB_2_4_port, Y => 
                           n947);
   U1318 : NAND3X1 port map( A => n945, B => n946, C => n947, Y => 
                           CARRYB_3_3_port);
   U1319 : XOR2X1 port map( A => n457, B => ab_6_3_port, Y => n948);
   U1320 : XOR2X1 port map( A => n526, B => n948, Y => SUMB_6_3_port);
   U1321 : NAND2X1 port map( A => SUMB_5_4_port, B => CARRYB_5_3_port, Y => 
                           n949);
   U1322 : NAND2X1 port map( A => SUMB_5_4_port, B => ab_6_3_port, Y => n950);
   U1323 : NAND2X1 port map( A => CARRYB_5_3_port, B => ab_6_3_port, Y => n951)
                           ;
   U1324 : NAND3X1 port map( A => n950, B => n949, C => n951, Y => 
                           CARRYB_6_3_port);
   U1325 : INVX2 port map( A => n999, Y => n973);
   U1326 : BUFX4 port map( A => CARRYB_2_0_port, Y => n968);
   U1327 : AND2X2 port map( A => SUMB_15_2_port, B => CARRYB_15_1_port, Y => 
                           n953);
   U1328 : AND2X2 port map( A => ab_0_1_port, B => ab_1_0_port, Y => n958);
   U1329 : AND2X2 port map( A => ab_0_4_port, B => ab_1_3_port, Y => n959);
   U1330 : AND2X2 port map( A => ab_0_3_port, B => ab_1_2_port, Y => n960);
   U1331 : NOR2X1 port map( A => n999, B => n655, Y => n962);
   U1332 : INVX2 port map( A => A(13), Y => n1054);
   U1333 : INVX2 port map( A => A(15), Y => n1052);
   U1334 : INVX2 port map( A => A(14), Y => n1053);
   U1335 : INVX2 port map( A => A(4), Y => n1023);
   U1336 : INVX2 port map( A => A(5), Y => n1025);
   U1337 : INVX2 port map( A => A(6), Y => n1027);
   U1338 : INVX2 port map( A => A(7), Y => n1029);
   U1339 : INVX2 port map( A => A(8), Y => n1031);
   U1340 : INVX2 port map( A => A(9), Y => n1033);
   U1341 : INVX2 port map( A => A(10), Y => n1035);
   U1342 : XOR2X1 port map( A => CARRYB_15_0_port, B => SUMB_15_1_port, Y => 
                           A1_14_port);
   U1343 : XOR2X1 port map( A => SUMB_15_2_port, B => CARRYB_15_1_port, Y => 
                           A1_15_port);
   U1344 : XOR2X1 port map( A => SUMB_15_4_port, B => CARRYB_15_3_port, Y => 
                           A1_17_port);
   U1345 : XOR2X1 port map( A => SUMB_15_6_port, B => CARRYB_15_5_port, Y => 
                           A1_19_port);
   U1346 : NAND2X1 port map( A => SUMB_15_7_port, B => CARRYB_15_6_port, Y => 
                           n963);
   U1347 : INVX2 port map( A => n963, Y => A2_21_port);
   U1348 : XOR2X1 port map( A => SUMB_15_8_port, B => CARRYB_15_7_port, Y => 
                           A1_21_port);
   U1349 : NAND2X1 port map( A => SUMB_15_8_port, B => CARRYB_15_7_port, Y => 
                           n964);
   U1350 : INVX2 port map( A => n964, Y => A2_22_port);
   U1351 : XOR2X1 port map( A => SUMB_15_9_port, B => CARRYB_15_8_port, Y => 
                           A1_22_port);
   U1352 : XOR2X1 port map( A => SUMB_15_10_port, B => CARRYB_15_9_port, Y => 
                           A1_23_port);
   U1353 : XOR2X1 port map( A => SUMB_15_11_port, B => CARRYB_15_10_port, Y => 
                           A1_24_port);
   U1354 : XOR2X1 port map( A => SUMB_15_12_port, B => CARRYB_15_11_port, Y => 
                           A1_25_port);
   U1355 : XOR2X1 port map( A => SUMB_15_13_port, B => CARRYB_15_12_port, Y => 
                           A1_26_port);
   U1356 : XOR2X1 port map( A => SUMB_15_14_port, B => CARRYB_15_13_port, Y => 
                           A1_27_port);
   U1357 : XOR2X1 port map( A => SUMB_15_15_port, B => CARRYB_15_14_port, Y => 
                           A1_28_port);
   U1358 : XOR2X1 port map( A => ab_1_0_port, B => ab_0_1_port, Y => PRODUCT(1)
                           );
   U1359 : XOR2X1 port map( A => ab_1_1_port, B => ab_0_2_port, Y => 
                           SUMB_1_1_port);
   U1360 : NAND2X1 port map( A => ab_0_2_port, B => ab_1_1_port, Y => n965);
   U1361 : INVX2 port map( A => n965, Y => CARRYB_1_1_port);
   U1362 : XOR2X1 port map( A => ab_1_2_port, B => ab_0_3_port, Y => 
                           SUMB_1_2_port);
   U1363 : XOR2X1 port map( A => ab_0_4_port, B => ab_1_3_port, Y => 
                           SUMB_1_3_port);
   U1364 : XOR2X1 port map( A => n962, B => ab_1_4_port, Y => SUMB_1_4_port);
   U1365 : XOR2X1 port map( A => ab_1_5_port, B => ab_0_6_port, Y => 
                           SUMB_1_5_port);
   U1366 : XOR2X1 port map( A => ab_1_6_port, B => ab_0_7_port, Y => 
                           SUMB_1_6_port);
   U1367 : XOR2X1 port map( A => ab_1_7_port, B => ab_0_8_port, Y => 
                           SUMB_1_7_port);
   U1368 : XOR2X1 port map( A => ab_1_8_port, B => ab_0_9_port, Y => 
                           SUMB_1_8_port);
   U1369 : XOR2X1 port map( A => ab_1_11_port, B => ab_0_12_port, Y => 
                           SUMB_1_11_port);
   U1370 : XOR2X1 port map( A => n96, B => ab_1_12_port, Y => SUMB_1_12_port);
   U1371 : NAND2X1 port map( A => ab_0_14_port, B => n139, Y => n966);
   U1372 : XOR2X1 port map( A => ab_1_14_port, B => n984, Y => SUMB_1_14_port);
   U1373 : BUFX4 port map( A => CARRYB_10_0_port, Y => n967);
   U1374 : INVX2 port map( A => n1000, Y => n1001);
   U1375 : INVX2 port map( A => B(6), Y => n1000);
   U1376 : INVX1 port map( A => n969, Y => n1044);
   U1377 : INVX2 port map( A => CARRYB_10_4_port, Y => n970);
   U1378 : INVX1 port map( A => n999, Y => n972);
   U1379 : INVX2 port map( A => B(5), Y => n999);
   U1380 : INVX2 port map( A => n989, Y => n990);
   U1381 : INVX1 port map( A => n973, Y => n1045);
   U1382 : INVX2 port map( A => CARRYB_2_4_port, Y => n975);
   U1383 : INVX2 port map( A => n993, Y => n976);
   U1384 : INVX2 port map( A => n993, Y => n994);
   U1385 : INVX2 port map( A => B(2), Y => n993);
   U1386 : INVX2 port map( A => n997, Y => n998);
   U1387 : INVX2 port map( A => n995, Y => n978);
   U1388 : INVX2 port map( A => n995, Y => n996);
   U1389 : INVX2 port map( A => B(3), Y => n995);
   U1390 : INVX1 port map( A => n977, Y => n1046);
   U1391 : INVX1 port map( A => n978, Y => n1047);
   U1392 : INVX2 port map( A => n991, Y => n992);
   U1393 : INVX2 port map( A => B(1), Y => n991);
   U1394 : INVX1 port map( A => n976, Y => n1048);
   U1395 : INVX1 port map( A => n980, Y => n1049);
   U1396 : INVX2 port map( A => n1016, Y => n985);
   U1397 : INVX2 port map( A => CARRYB_11_1_port, Y => n981);
   U1398 : INVX2 port map( A => CARRYB_2_3_port, Y => n983);
   U1399 : INVX4 port map( A => A(1), Y => n1017);
   U1400 : INVX2 port map( A => CARRYB_2_2_port, Y => n986);
   U1401 : INVX8 port map( A => n1014, Y => n1015);
   U1402 : INVX8 port map( A => n1021, Y => n1022);
   U1403 : INVX8 port map( A => n1023, Y => n1024);
   U1404 : INVX8 port map( A => n1025, Y => n1026);
   U1405 : INVX8 port map( A => n1027, Y => n1028);
   U1406 : INVX8 port map( A => n1029, Y => n1030);
   U1407 : INVX8 port map( A => n1031, Y => n1032);
   U1408 : INVX8 port map( A => n1033, Y => n1034);
   U1409 : INVX8 port map( A => n1035, Y => n1036);
   U1410 : AND2X2 port map( A => n1018, B => B(14), Y => ab_1_14_port);
   U1411 : AND2X2 port map( A => B(14), B => n401, Y => ab_0_14_port);
   U1412 : AND2X2 port map( A => n1018, B => B(12), Y => ab_1_12_port);
   U1413 : AND2X2 port map( A => B(12), B => n531, Y => ab_0_12_port);
   U1414 : AND2X2 port map( A => n423, B => B(10), Y => ab_1_10_port);
   U1415 : AND2X2 port map( A => n531, B => B(10), Y => ab_0_10_port);
   U1416 : AND2X2 port map( A => B(9), B => n531, Y => ab_0_9_port);
   U1417 : AND2X2 port map( A => n1018, B => B(8), Y => ab_1_8_port);
   U1418 : AND2X2 port map( A => n985, B => B(8), Y => ab_0_8_port);
   U1419 : AND2X2 port map( A => n1003, B => n423, Y => ab_1_7_port);
   U1420 : AND2X2 port map( A => n1003, B => n985, Y => ab_0_7_port);
   U1421 : AND2X2 port map( A => n1018, B => n1001, Y => ab_1_6_port);
   U1422 : AND2X2 port map( A => n1001, B => n402, Y => ab_0_6_port);
   U1423 : AND2X2 port map( A => B(5), B => n1018, Y => ab_1_5_port);
   U1424 : AND2X2 port map( A => n1018, B => n998, Y => ab_1_4_port);
   U1425 : AND2X2 port map( A => n998, B => n402, Y => ab_0_4_port);
   U1426 : AND2X2 port map( A => n1018, B => n996, Y => ab_1_3_port);
   U1427 : AND2X2 port map( A => n996, B => n401, Y => ab_0_3_port);
   U1428 : AND2X2 port map( A => n994, B => n9, Y => ab_1_2_port);
   U1429 : AND2X2 port map( A => n994, B => n402, Y => ab_0_2_port);
   U1430 : AND2X2 port map( A => n1018, B => n992, Y => ab_1_1_port);
   U1431 : AND2X2 port map( A => n992, B => n402, Y => ab_0_1_port);
   U1432 : AND2X2 port map( A => n9, B => n990, Y => ab_1_0_port);
   U1433 : NOR2X1 port map( A => n1018, B => n1051, Y => ab_1_15_port);
   U1434 : AND2X2 port map( A => n4, B => n1013, Y => ab_2_13_port);
   U1435 : AND2X2 port map( A => n5, B => n1011, Y => ab_2_12_port);
   U1436 : AND2X2 port map( A => n5, B => n1009, Y => ab_2_11_port);
   U1437 : AND2X2 port map( A => n1020, B => n1007, Y => ab_2_10_port);
   U1438 : AND2X2 port map( A => n1020, B => B(9), Y => ab_2_9_port);
   U1439 : AND2X2 port map( A => n1020, B => B(8), Y => ab_2_8_port);
   U1440 : AND2X2 port map( A => n4, B => n969, Y => ab_2_6_port);
   U1441 : AND2X2 port map( A => n5, B => n973, Y => ab_2_5_port);
   U1442 : AND2X2 port map( A => n4, B => n977, Y => ab_2_4_port);
   U1443 : AND2X2 port map( A => n10, B => n978, Y => ab_2_3_port);
   U1444 : AND2X2 port map( A => n10, B => n976, Y => ab_2_2_port);
   U1445 : AND2X2 port map( A => n5, B => n980, Y => ab_2_1_port);
   U1446 : AND2X2 port map( A => n5, B => n974, Y => ab_2_0_port);
   U1447 : AND2X2 port map( A => n1022, B => n1015, Y => ab_3_14_port);
   U1448 : NOR2X1 port map( A => n4, B => n1051, Y => ab_2_15_port);
   U1449 : AND2X2 port map( A => n1022, B => n1013, Y => ab_3_13_port);
   U1450 : AND2X2 port map( A => n1022, B => n1011, Y => ab_3_12_port);
   U1451 : AND2X2 port map( A => n1022, B => n1009, Y => ab_3_11_port);
   U1452 : AND2X2 port map( A => n1022, B => n1007, Y => ab_3_10_port);
   U1453 : AND2X2 port map( A => n1022, B => n507, Y => ab_3_9_port);
   U1454 : AND2X2 port map( A => n1022, B => n905, Y => ab_3_7_port);
   U1455 : AND2X2 port map( A => n1022, B => n969, Y => ab_3_6_port);
   U1456 : AND2X2 port map( A => n1022, B => n972, Y => ab_3_5_port);
   U1457 : AND2X2 port map( A => n1022, B => n977, Y => ab_3_4_port);
   U1458 : AND2X2 port map( A => n1022, B => n978, Y => ab_3_3_port);
   U1459 : AND2X2 port map( A => n1022, B => n976, Y => ab_3_2_port);
   U1460 : AND2X2 port map( A => n1022, B => n980, Y => ab_3_1_port);
   U1461 : AND2X2 port map( A => n1022, B => n974, Y => ab_3_0_port);
   U1462 : AND2X2 port map( A => n1024, B => n1015, Y => ab_4_14_port);
   U1463 : NOR2X1 port map( A => n1022, B => n1051, Y => ab_3_15_port);
   U1464 : AND2X2 port map( A => n1024, B => n1013, Y => ab_4_13_port);
   U1465 : AND2X2 port map( A => n1024, B => n1011, Y => ab_4_12_port);
   U1466 : AND2X2 port map( A => n1024, B => n1009, Y => ab_4_11_port);
   U1467 : AND2X2 port map( A => n1024, B => n1007, Y => ab_4_10_port);
   U1468 : AND2X2 port map( A => n1024, B => n507, Y => ab_4_9_port);
   U1469 : AND2X2 port map( A => n1024, B => n1005, Y => ab_4_8_port);
   U1470 : AND2X2 port map( A => n1024, B => n905, Y => ab_4_7_port);
   U1471 : AND2X2 port map( A => n1024, B => n969, Y => ab_4_6_port);
   U1472 : AND2X2 port map( A => n1024, B => n973, Y => ab_4_5_port);
   U1473 : AND2X2 port map( A => n1024, B => n977, Y => ab_4_4_port);
   U1474 : AND2X2 port map( A => n1024, B => n978, Y => ab_4_3_port);
   U1475 : AND2X2 port map( A => n1024, B => n976, Y => ab_4_2_port);
   U1476 : AND2X2 port map( A => n1024, B => n980, Y => ab_4_1_port);
   U1477 : AND2X2 port map( A => n1024, B => n974, Y => ab_4_0_port);
   U1478 : AND2X2 port map( A => n1026, B => n1015, Y => ab_5_14_port);
   U1479 : NOR2X1 port map( A => n1024, B => n1051, Y => ab_4_15_port);
   U1480 : AND2X2 port map( A => n1026, B => n1013, Y => ab_5_13_port);
   U1481 : AND2X2 port map( A => n1026, B => n1011, Y => ab_5_12_port);
   U1482 : AND2X2 port map( A => n1026, B => n163, Y => ab_5_11_port);
   U1483 : AND2X2 port map( A => n1026, B => n1007, Y => ab_5_10_port);
   U1484 : AND2X2 port map( A => n1026, B => n507, Y => ab_5_9_port);
   U1485 : AND2X2 port map( A => n1026, B => n1005, Y => ab_5_8_port);
   U1486 : AND2X2 port map( A => n1026, B => n905, Y => ab_5_7_port);
   U1487 : AND2X2 port map( A => n1026, B => n969, Y => ab_5_6_port);
   U1488 : AND2X2 port map( A => n1026, B => n972, Y => ab_5_5_port);
   U1489 : AND2X2 port map( A => n1026, B => n977, Y => ab_5_4_port);
   U1490 : AND2X2 port map( A => n1026, B => n978, Y => ab_5_3_port);
   U1491 : AND2X2 port map( A => n1026, B => n976, Y => ab_5_2_port);
   U1492 : AND2X2 port map( A => n1026, B => n980, Y => ab_5_1_port);
   U1493 : AND2X2 port map( A => n1026, B => n974, Y => ab_5_0_port);
   U1494 : AND2X2 port map( A => n1028, B => n1015, Y => ab_6_14_port);
   U1495 : NOR2X1 port map( A => n1026, B => n1051, Y => ab_5_15_port);
   U1496 : AND2X2 port map( A => n1028, B => n1013, Y => ab_6_13_port);
   U1497 : AND2X2 port map( A => n1028, B => n1011, Y => ab_6_12_port);
   U1498 : AND2X2 port map( A => n1028, B => n163, Y => ab_6_11_port);
   U1499 : AND2X2 port map( A => n1028, B => n1007, Y => ab_6_10_port);
   U1500 : AND2X2 port map( A => n1028, B => n507, Y => ab_6_9_port);
   U1501 : AND2X2 port map( A => n1028, B => n1005, Y => ab_6_8_port);
   U1502 : AND2X2 port map( A => n1028, B => n905, Y => ab_6_7_port);
   U1503 : AND2X2 port map( A => n1028, B => n969, Y => ab_6_6_port);
   U1504 : AND2X2 port map( A => n1028, B => n973, Y => ab_6_5_port);
   U1505 : AND2X2 port map( A => n1028, B => n977, Y => ab_6_4_port);
   U1506 : AND2X2 port map( A => n1028, B => n978, Y => ab_6_3_port);
   U1507 : AND2X2 port map( A => n1028, B => n976, Y => ab_6_2_port);
   U1508 : AND2X2 port map( A => n1028, B => n980, Y => ab_6_1_port);
   U1509 : AND2X2 port map( A => n1028, B => n974, Y => ab_6_0_port);
   U1510 : AND2X2 port map( A => n1030, B => n1015, Y => ab_7_14_port);
   U1511 : NOR2X1 port map( A => n1028, B => n1051, Y => ab_6_15_port);
   U1512 : AND2X2 port map( A => n1030, B => n1013, Y => ab_7_13_port);
   U1513 : AND2X2 port map( A => n1030, B => n1011, Y => ab_7_12_port);
   U1514 : AND2X2 port map( A => n1030, B => n163, Y => ab_7_11_port);
   U1515 : AND2X2 port map( A => n1030, B => n1007, Y => ab_7_10_port);
   U1516 : AND2X2 port map( A => n1030, B => n507, Y => ab_7_9_port);
   U1517 : AND2X2 port map( A => n1030, B => n1005, Y => ab_7_8_port);
   U1518 : AND2X2 port map( A => n1030, B => n905, Y => ab_7_7_port);
   U1519 : AND2X2 port map( A => n1030, B => n969, Y => ab_7_6_port);
   U1520 : AND2X2 port map( A => n1030, B => n972, Y => ab_7_5_port);
   U1521 : AND2X2 port map( A => n1030, B => n977, Y => ab_7_4_port);
   U1522 : AND2X2 port map( A => n1030, B => n978, Y => ab_7_3_port);
   U1523 : AND2X2 port map( A => n1030, B => n976, Y => ab_7_2_port);
   U1524 : AND2X2 port map( A => n1030, B => n980, Y => ab_7_1_port);
   U1525 : AND2X2 port map( A => n1030, B => n974, Y => ab_7_0_port);
   U1526 : AND2X2 port map( A => n1032, B => n1015, Y => ab_8_14_port);
   U1527 : NOR2X1 port map( A => n1030, B => n1051, Y => ab_7_15_port);
   U1528 : AND2X2 port map( A => n1032, B => n1013, Y => ab_8_13_port);
   U1529 : AND2X2 port map( A => n1032, B => n1011, Y => ab_8_12_port);
   U1530 : AND2X2 port map( A => n1032, B => n163, Y => ab_8_11_port);
   U1531 : AND2X2 port map( A => n1032, B => n1007, Y => ab_8_10_port);
   U1532 : AND2X2 port map( A => n1032, B => n507, Y => ab_8_9_port);
   U1533 : AND2X2 port map( A => n1032, B => n1005, Y => ab_8_8_port);
   U1534 : AND2X2 port map( A => n1032, B => n905, Y => ab_8_7_port);
   U1535 : AND2X2 port map( A => n1032, B => n969, Y => ab_8_6_port);
   U1536 : AND2X2 port map( A => n1032, B => n973, Y => ab_8_5_port);
   U1537 : AND2X2 port map( A => n1032, B => n977, Y => ab_8_4_port);
   U1538 : AND2X2 port map( A => n1032, B => n978, Y => ab_8_3_port);
   U1539 : AND2X2 port map( A => n1032, B => n976, Y => ab_8_2_port);
   U1540 : AND2X2 port map( A => n1032, B => n980, Y => ab_8_1_port);
   U1541 : AND2X2 port map( A => n1032, B => n974, Y => ab_8_0_port);
   U1542 : AND2X2 port map( A => n1034, B => n1015, Y => ab_9_14_port);
   U1543 : NOR2X1 port map( A => n1032, B => n1051, Y => ab_8_15_port);
   U1544 : AND2X2 port map( A => n1034, B => n1013, Y => ab_9_13_port);
   U1545 : AND2X2 port map( A => n1034, B => n1011, Y => ab_9_12_port);
   U1546 : AND2X2 port map( A => n1034, B => n163, Y => ab_9_11_port);
   U1547 : AND2X2 port map( A => n1034, B => n1007, Y => ab_9_10_port);
   U1548 : AND2X2 port map( A => n1034, B => n507, Y => ab_9_9_port);
   U1549 : AND2X2 port map( A => n1034, B => n1005, Y => ab_9_8_port);
   U1550 : AND2X2 port map( A => n1034, B => n905, Y => ab_9_7_port);
   U1551 : AND2X2 port map( A => n1034, B => n969, Y => ab_9_6_port);
   U1552 : AND2X2 port map( A => n1034, B => n972, Y => ab_9_5_port);
   U1553 : AND2X2 port map( A => n1034, B => n977, Y => ab_9_4_port);
   U1554 : AND2X2 port map( A => n1034, B => n978, Y => ab_9_3_port);
   U1555 : AND2X2 port map( A => n1034, B => n976, Y => ab_9_2_port);
   U1556 : AND2X2 port map( A => n1034, B => n980, Y => ab_9_1_port);
   U1557 : AND2X2 port map( A => n1034, B => n974, Y => ab_9_0_port);
   U1558 : AND2X2 port map( A => n1036, B => n1015, Y => ab_10_14_port);
   U1559 : NOR2X1 port map( A => n1034, B => n1051, Y => ab_9_15_port);
   U1560 : AND2X2 port map( A => n1036, B => n1013, Y => ab_10_13_port);
   U1561 : AND2X2 port map( A => n1036, B => n1011, Y => ab_10_12_port);
   U1562 : AND2X2 port map( A => n1036, B => n163, Y => ab_10_11_port);
   U1563 : AND2X2 port map( A => n1036, B => n1007, Y => ab_10_10_port);
   U1564 : AND2X2 port map( A => n1036, B => n507, Y => ab_10_9_port);
   U1565 : AND2X2 port map( A => n1036, B => n1005, Y => ab_10_8_port);
   U1566 : AND2X2 port map( A => n1036, B => n905, Y => ab_10_7_port);
   U1567 : AND2X2 port map( A => n1036, B => n969, Y => ab_10_6_port);
   U1568 : AND2X2 port map( A => n1036, B => n973, Y => ab_10_5_port);
   U1569 : AND2X2 port map( A => n1036, B => n977, Y => ab_10_4_port);
   U1570 : AND2X2 port map( A => n1036, B => n978, Y => ab_10_3_port);
   U1571 : AND2X2 port map( A => n1036, B => n976, Y => ab_10_2_port);
   U1572 : AND2X2 port map( A => n1036, B => n980, Y => ab_10_1_port);
   U1573 : AND2X2 port map( A => n1036, B => n974, Y => ab_10_0_port);
   U1574 : AND2X2 port map( A => A(11), B => n1015, Y => ab_11_14_port);
   U1575 : NOR2X1 port map( A => n1036, B => n1051, Y => ab_10_15_port);
   U1576 : AND2X2 port map( A => A(11), B => n1013, Y => ab_11_13_port);
   U1577 : AND2X2 port map( A => A(11), B => n1011, Y => ab_11_12_port);
   U1578 : AND2X2 port map( A => A(11), B => n163, Y => ab_11_11_port);
   U1579 : AND2X2 port map( A => A(11), B => n1007, Y => ab_11_10_port);
   U1580 : AND2X2 port map( A => A(11), B => n507, Y => ab_11_9_port);
   U1581 : AND2X2 port map( A => A(11), B => n1005, Y => ab_11_8_port);
   U1582 : AND2X2 port map( A => A(11), B => n905, Y => ab_11_7_port);
   U1583 : AND2X2 port map( A => A(11), B => n969, Y => ab_11_6_port);
   U1584 : AND2X2 port map( A => A(11), B => n972, Y => ab_11_5_port);
   U1585 : AND2X2 port map( A => A(11), B => n977, Y => ab_11_4_port);
   U1586 : AND2X2 port map( A => A(11), B => n978, Y => ab_11_3_port);
   U1587 : AND2X2 port map( A => A(11), B => n976, Y => ab_11_2_port);
   U1588 : AND2X2 port map( A => A(11), B => n980, Y => ab_11_1_port);
   U1589 : AND2X2 port map( A => A(11), B => n974, Y => ab_11_0_port);
   U1590 : AND2X2 port map( A => A(12), B => n1015, Y => ab_12_14_port);
   U1591 : NOR2X1 port map( A => A(11), B => n1051, Y => ab_11_15_port);
   U1592 : AND2X2 port map( A => A(12), B => n1013, Y => ab_12_13_port);
   U1593 : AND2X2 port map( A => A(12), B => n1011, Y => ab_12_12_port);
   U1594 : AND2X2 port map( A => A(12), B => n163, Y => ab_12_11_port);
   U1595 : AND2X2 port map( A => A(12), B => n1007, Y => ab_12_10_port);
   U1596 : AND2X2 port map( A => A(12), B => n507, Y => ab_12_9_port);
   U1597 : AND2X2 port map( A => A(12), B => n1005, Y => ab_12_8_port);
   U1598 : AND2X2 port map( A => A(12), B => n905, Y => ab_12_7_port);
   U1599 : AND2X2 port map( A => A(12), B => n969, Y => ab_12_6_port);
   U1600 : AND2X2 port map( A => A(12), B => n973, Y => ab_12_5_port);
   U1601 : AND2X2 port map( A => A(12), B => n977, Y => ab_12_4_port);
   U1602 : AND2X2 port map( A => A(12), B => n978, Y => ab_12_3_port);
   U1603 : AND2X2 port map( A => A(12), B => n976, Y => ab_12_2_port);
   U1604 : AND2X2 port map( A => A(12), B => n980, Y => ab_12_1_port);
   U1605 : AND2X2 port map( A => A(12), B => n974, Y => ab_12_0_port);
   U1606 : NOR2X1 port map( A => n1054, B => n1037, Y => ab_13_14_port);
   U1607 : NOR2X1 port map( A => A(12), B => n1051, Y => ab_12_15_port);
   U1608 : NOR2X1 port map( A => n1054, B => n1038, Y => ab_13_13_port);
   U1609 : NOR2X1 port map( A => n1054, B => n1039, Y => ab_13_12_port);
   U1610 : NOR2X1 port map( A => n1054, B => n1040, Y => ab_13_11_port);
   U1611 : NOR2X1 port map( A => n1054, B => n1041, Y => ab_13_10_port);
   U1612 : NOR2X1 port map( A => n1054, B => n1042, Y => ab_13_9_port);
   U1613 : NOR2X1 port map( A => n1054, B => n1004, Y => ab_13_8_port);
   U1614 : NOR2X1 port map( A => n1054, B => n1043, Y => ab_13_7_port);
   U1615 : NOR2X1 port map( A => n1054, B => n1044, Y => ab_13_6_port);
   U1616 : NOR2X1 port map( A => n1054, B => n1045, Y => ab_13_5_port);
   U1617 : NOR2X1 port map( A => n1054, B => n1046, Y => ab_13_4_port);
   U1618 : NOR2X1 port map( A => n1054, B => n1047, Y => ab_13_3_port);
   U1619 : NOR2X1 port map( A => n1054, B => n1048, Y => ab_13_2_port);
   U1620 : NOR2X1 port map( A => n1054, B => n1049, Y => ab_13_1_port);
   U1621 : NOR2X1 port map( A => n1054, B => n989, Y => ab_13_0_port);
   U1622 : NOR2X1 port map( A => n1053, B => n1037, Y => ab_14_14_port);
   U1623 : NOR2X1 port map( A => A(13), B => n1051, Y => ab_13_15_port);
   U1624 : NOR2X1 port map( A => n1053, B => n1038, Y => ab_14_13_port);
   U1625 : NOR2X1 port map( A => n1053, B => n1039, Y => ab_14_12_port);
   U1626 : NOR2X1 port map( A => n1053, B => n1040, Y => ab_14_11_port);
   U1627 : NOR2X1 port map( A => n1053, B => n1041, Y => ab_14_10_port);
   U1628 : NOR2X1 port map( A => n1053, B => n1042, Y => ab_14_9_port);
   U1629 : NOR2X1 port map( A => n1053, B => n1004, Y => ab_14_8_port);
   U1630 : NOR2X1 port map( A => n1053, B => n1043, Y => ab_14_7_port);
   U1631 : NOR2X1 port map( A => n1053, B => n1044, Y => ab_14_6_port);
   U1632 : NOR2X1 port map( A => n1053, B => n1045, Y => ab_14_5_port);
   U1633 : NOR2X1 port map( A => n1053, B => n1046, Y => ab_14_4_port);
   U1634 : NOR2X1 port map( A => n1053, B => n1047, Y => ab_14_3_port);
   U1635 : NOR2X1 port map( A => n1053, B => n1048, Y => ab_14_2_port);
   U1636 : NOR2X1 port map( A => n1053, B => n1049, Y => ab_14_1_port);
   U1637 : NOR2X1 port map( A => n1053, B => n989, Y => ab_14_0_port);
   U1638 : NOR2X1 port map( A => n1052, B => n1051, Y => ab_15_15_port);
   U1639 : NOR2X1 port map( A => A(14), B => n1051, Y => ab_14_15_port);
   U1640 : AND2X2 port map( A => n974, B => n402, Y => PRODUCT(0));
   U1641 : INVX2 port map( A => CARRYB_15_15_port, Y => n1050);
   U1642 : NOR2X1 port map( A => n507, B => n1052, Y => ab_15_9_port);
   U1643 : NOR2X1 port map( A => n1005, B => n1052, Y => ab_15_8_port);
   U1644 : NOR2X1 port map( A => n905, B => n1052, Y => ab_15_7_port);
   U1645 : NOR2X1 port map( A => n969, B => n1052, Y => ab_15_6_port);
   U1646 : NOR2X1 port map( A => n972, B => n1052, Y => ab_15_5_port);
   U1647 : NOR2X1 port map( A => n977, B => n1052, Y => ab_15_4_port);
   U1648 : NOR2X1 port map( A => n978, B => n1052, Y => ab_15_3_port);
   U1649 : NOR2X1 port map( A => n976, B => n1052, Y => ab_15_2_port);
   U1650 : NOR2X1 port map( A => n980, B => n1052, Y => ab_15_1_port);
   U1651 : NOR2X1 port map( A => n1015, B => n1052, Y => ab_15_14_port);
   U1652 : NOR2X1 port map( A => n1013, B => n1052, Y => ab_15_13_port);
   U1653 : NOR2X1 port map( A => n1011, B => n1052, Y => ab_15_12_port);
   U1654 : NOR2X1 port map( A => n163, B => n1052, Y => ab_15_11_port);
   U1655 : NOR2X1 port map( A => n1007, B => n1052, Y => ab_15_10_port);
   U1656 : NOR2X1 port map( A => n974, B => n1052, Y => ab_15_0_port);
   n1055 <= '0';

end SYN_csa;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW02_mult_1 is

   port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  PRODUCT
         : out std_logic_vector (31 downto 0));

end matrix_math_DW02_mult_1;

architecture SYN_csa of matrix_math_DW02_mult_1 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component matrix_math_DW01_add_23
      port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (29 downto 0);  CO : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_15_15_port, ab_15_14_port, ab_15_13_port, 
      ab_15_12_port, ab_15_11_port, ab_15_10_port, ab_15_9_port, ab_15_8_port, 
      ab_15_7_port, ab_15_6_port, ab_15_5_port, ab_15_4_port, ab_15_3_port, 
      ab_15_2_port, ab_15_1_port, ab_15_0_port, ab_14_15_port, ab_14_14_port, 
      ab_14_13_port, ab_14_12_port, ab_14_11_port, ab_14_10_port, ab_14_9_port,
      ab_14_8_port, ab_14_7_port, ab_14_6_port, ab_14_5_port, ab_14_4_port, 
      ab_14_3_port, ab_14_2_port, ab_14_1_port, ab_14_0_port, ab_13_15_port, 
      ab_13_14_port, ab_13_13_port, ab_13_12_port, ab_13_11_port, ab_13_10_port
      , ab_13_9_port, ab_13_8_port, ab_13_7_port, ab_13_6_port, ab_13_5_port, 
      ab_13_4_port, ab_13_3_port, ab_13_2_port, ab_13_1_port, ab_13_0_port, 
      ab_12_15_port, ab_12_14_port, ab_12_13_port, ab_12_12_port, ab_12_11_port
      , ab_12_10_port, ab_12_9_port, ab_12_8_port, ab_12_7_port, ab_12_6_port, 
      ab_12_5_port, ab_12_4_port, ab_12_3_port, ab_12_2_port, ab_12_1_port, 
      ab_12_0_port, ab_11_15_port, ab_11_14_port, ab_11_13_port, ab_11_12_port,
      ab_11_11_port, ab_11_10_port, ab_11_9_port, ab_11_8_port, ab_11_7_port, 
      ab_11_6_port, ab_11_5_port, ab_11_4_port, ab_11_3_port, ab_11_2_port, 
      ab_11_1_port, ab_11_0_port, ab_10_15_port, ab_10_14_port, ab_10_13_port, 
      ab_10_12_port, ab_10_11_port, ab_10_10_port, ab_10_9_port, ab_10_8_port, 
      ab_10_7_port, ab_10_6_port, ab_10_5_port, ab_10_4_port, ab_10_3_port, 
      ab_10_2_port, ab_10_1_port, ab_10_0_port, ab_9_15_port, ab_9_14_port, 
      ab_9_13_port, ab_9_12_port, ab_9_11_port, ab_9_10_port, ab_9_9_port, 
      ab_9_8_port, ab_9_7_port, ab_9_6_port, ab_9_5_port, ab_9_4_port, 
      ab_9_3_port, ab_9_2_port, ab_9_1_port, ab_9_0_port, ab_8_15_port, 
      ab_8_14_port, ab_8_13_port, ab_8_12_port, ab_8_11_port, ab_8_10_port, 
      ab_8_9_port, ab_8_8_port, ab_8_7_port, ab_8_6_port, ab_8_5_port, 
      ab_8_4_port, ab_8_3_port, ab_8_2_port, ab_8_1_port, ab_8_0_port, 
      ab_7_15_port, ab_7_14_port, ab_7_13_port, ab_7_12_port, ab_7_11_port, 
      ab_7_10_port, ab_7_9_port, ab_7_8_port, ab_7_7_port, ab_7_6_port, 
      ab_7_5_port, ab_7_4_port, ab_7_3_port, ab_7_2_port, ab_7_1_port, 
      ab_7_0_port, ab_6_15_port, ab_6_14_port, ab_6_13_port, ab_6_12_port, 
      ab_6_11_port, ab_6_10_port, ab_6_9_port, ab_6_8_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_15_port, ab_5_14_port, ab_5_13_port, 
      ab_5_12_port, ab_5_11_port, ab_5_10_port, ab_5_9_port, ab_5_8_port, 
      ab_5_7_port, ab_5_6_port, ab_5_5_port, ab_5_4_port, ab_5_3_port, 
      ab_5_2_port, ab_5_1_port, ab_5_0_port, ab_4_15_port, ab_4_14_port, 
      ab_4_13_port, ab_4_12_port, ab_4_11_port, ab_4_10_port, ab_4_9_port, 
      ab_4_8_port, ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, 
      ab_4_3_port, ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_15_port, 
      ab_3_14_port, ab_3_13_port, ab_3_12_port, ab_3_11_port, ab_3_10_port, 
      ab_3_9_port, ab_3_8_port, ab_3_7_port, ab_3_6_port, ab_3_5_port, 
      ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, ab_3_0_port, 
      ab_2_15_port, ab_2_14_port, ab_2_13_port, ab_2_12_port, ab_2_11_port, 
      ab_2_10_port, ab_2_9_port, ab_2_8_port, ab_2_7_port, ab_2_6_port, 
      ab_2_5_port, ab_2_4_port, ab_2_3_port, ab_2_2_port, ab_2_1_port, 
      ab_2_0_port, ab_1_15_port, ab_1_14_port, ab_1_13_port, ab_1_12_port, 
      ab_1_11_port, ab_1_10_port, ab_1_8_port, ab_1_7_port, ab_1_6_port, 
      ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_1_port, ab_1_0_port, 
      ab_0_15_port, ab_0_14_port, ab_0_13_port, ab_0_12_port, ab_0_11_port, 
      ab_0_10_port, ab_0_9_port, ab_0_8_port, ab_0_7_port, ab_0_6_port, 
      ab_0_5_port, ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, 
      CARRYB_15_15_port, CARRYB_15_14_port, CARRYB_15_13_port, 
      CARRYB_15_12_port, CARRYB_15_11_port, CARRYB_15_10_port, CARRYB_15_9_port
      , CARRYB_15_8_port, CARRYB_15_7_port, CARRYB_15_6_port, CARRYB_15_5_port,
      CARRYB_15_4_port, CARRYB_15_3_port, CARRYB_15_2_port, CARRYB_15_1_port, 
      CARRYB_15_0_port, CARRYB_14_14_port, CARRYB_14_13_port, CARRYB_14_12_port
      , CARRYB_14_11_port, CARRYB_14_10_port, CARRYB_14_9_port, 
      CARRYB_14_8_port, CARRYB_14_7_port, CARRYB_14_6_port, CARRYB_14_5_port, 
      CARRYB_14_4_port, CARRYB_14_3_port, CARRYB_14_2_port, CARRYB_14_1_port, 
      CARRYB_14_0_port, CARRYB_13_14_port, CARRYB_13_13_port, CARRYB_13_12_port
      , CARRYB_13_11_port, CARRYB_13_10_port, CARRYB_13_9_port, 
      CARRYB_13_8_port, CARRYB_13_7_port, CARRYB_13_6_port, CARRYB_13_5_port, 
      CARRYB_13_4_port, CARRYB_13_3_port, CARRYB_13_2_port, CARRYB_13_1_port, 
      CARRYB_13_0_port, CARRYB_12_14_port, CARRYB_12_13_port, CARRYB_12_12_port
      , CARRYB_12_11_port, CARRYB_12_10_port, CARRYB_12_9_port, 
      CARRYB_12_8_port, CARRYB_12_7_port, CARRYB_12_6_port, CARRYB_12_5_port, 
      CARRYB_12_4_port, CARRYB_12_3_port, CARRYB_12_2_port, CARRYB_12_1_port, 
      CARRYB_12_0_port, CARRYB_11_14_port, CARRYB_11_13_port, CARRYB_11_12_port
      , CARRYB_11_11_port, CARRYB_11_10_port, CARRYB_11_9_port, 
      CARRYB_11_8_port, CARRYB_11_7_port, CARRYB_11_6_port, CARRYB_11_5_port, 
      CARRYB_11_4_port, CARRYB_11_3_port, CARRYB_11_2_port, CARRYB_11_1_port, 
      CARRYB_11_0_port, CARRYB_10_14_port, CARRYB_10_13_port, CARRYB_10_12_port
      , CARRYB_10_11_port, CARRYB_10_10_port, CARRYB_10_9_port, 
      CARRYB_10_8_port, CARRYB_10_7_port, CARRYB_10_6_port, CARRYB_10_5_port, 
      CARRYB_10_4_port, CARRYB_10_3_port, CARRYB_10_1_port, CARRYB_10_0_port, 
      CARRYB_9_14_port, CARRYB_9_13_port, CARRYB_9_12_port, CARRYB_9_11_port, 
      CARRYB_9_10_port, CARRYB_9_9_port, CARRYB_9_8_port, CARRYB_9_7_port, 
      CARRYB_9_6_port, CARRYB_9_5_port, CARRYB_9_4_port, CARRYB_9_3_port, 
      CARRYB_9_2_port, CARRYB_9_1_port, CARRYB_9_0_port, CARRYB_8_14_port, 
      CARRYB_8_13_port, CARRYB_8_12_port, CARRYB_8_11_port, CARRYB_8_10_port, 
      CARRYB_8_9_port, CARRYB_8_8_port, CARRYB_8_7_port, CARRYB_8_6_port, 
      CARRYB_8_5_port, CARRYB_8_4_port, CARRYB_8_3_port, CARRYB_8_2_port, 
      CARRYB_8_1_port, CARRYB_8_0_port, CARRYB_7_14_port, CARRYB_7_13_port, 
      CARRYB_7_12_port, CARRYB_7_11_port, CARRYB_7_10_port, CARRYB_7_9_port, 
      CARRYB_7_8_port, CARRYB_7_7_port, CARRYB_7_6_port, CARRYB_7_5_port, 
      CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, CARRYB_7_1_port, 
      CARRYB_7_0_port, CARRYB_6_14_port, CARRYB_6_13_port, CARRYB_6_12_port, 
      CARRYB_6_11_port, CARRYB_6_10_port, CARRYB_6_9_port, CARRYB_6_8_port, 
      CARRYB_6_7_port, CARRYB_6_6_port, CARRYB_6_5_port, CARRYB_6_4_port, 
      CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, CARRYB_6_0_port, 
      CARRYB_5_14_port, CARRYB_5_13_port, CARRYB_5_12_port, CARRYB_5_11_port, 
      CARRYB_5_10_port, CARRYB_5_9_port, CARRYB_5_8_port, CARRYB_5_7_port, 
      CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, CARRYB_5_2_port, 
      CARRYB_5_1_port, CARRYB_5_0_port, CARRYB_4_14_port, CARRYB_4_13_port, 
      CARRYB_4_12_port, CARRYB_4_11_port, CARRYB_4_10_port, CARRYB_4_9_port, 
      CARRYB_4_8_port, CARRYB_4_7_port, CARRYB_4_6_port, CARRYB_4_5_port, 
      CARRYB_4_4_port, CARRYB_4_3_port, CARRYB_4_2_port, CARRYB_4_1_port, 
      CARRYB_4_0_port, CARRYB_3_14_port, CARRYB_3_13_port, CARRYB_3_12_port, 
      CARRYB_3_11_port, CARRYB_3_10_port, CARRYB_3_9_port, CARRYB_3_8_port, 
      CARRYB_3_7_port, CARRYB_3_6_port, CARRYB_3_5_port, CARRYB_3_4_port, 
      CARRYB_3_3_port, CARRYB_3_2_port, CARRYB_3_1_port, CARRYB_3_0_port, 
      CARRYB_2_14_port, CARRYB_2_13_port, CARRYB_2_12_port, CARRYB_2_11_port, 
      CARRYB_2_10_port, CARRYB_2_9_port, CARRYB_2_8_port, CARRYB_2_7_port, 
      CARRYB_2_6_port, CARRYB_2_5_port, CARRYB_2_4_port, CARRYB_2_3_port, 
      CARRYB_2_2_port, CARRYB_2_1_port, CARRYB_2_0_port, CARRYB_1_13_port, 
      SUMB_15_15_port, SUMB_15_14_port, SUMB_15_13_port, SUMB_15_12_port, 
      SUMB_15_11_port, SUMB_15_10_port, SUMB_15_9_port, SUMB_15_8_port, 
      SUMB_15_7_port, SUMB_15_6_port, SUMB_15_5_port, SUMB_15_4_port, 
      SUMB_15_3_port, SUMB_15_2_port, SUMB_15_1_port, SUMB_15_0_port, 
      SUMB_14_14_port, SUMB_14_13_port, SUMB_14_12_port, SUMB_14_11_port, 
      SUMB_14_10_port, SUMB_14_9_port, SUMB_14_8_port, SUMB_14_7_port, 
      SUMB_14_6_port, SUMB_14_5_port, SUMB_14_4_port, SUMB_14_3_port, 
      SUMB_14_2_port, SUMB_14_1_port, SUMB_13_14_port, SUMB_13_13_port, 
      SUMB_13_12_port, SUMB_13_11_port, SUMB_13_10_port, SUMB_13_9_port, 
      SUMB_13_8_port, SUMB_13_7_port, SUMB_13_6_port, SUMB_13_5_port, 
      SUMB_13_4_port, SUMB_13_3_port, SUMB_13_2_port, SUMB_13_1_port, 
      SUMB_12_14_port, SUMB_12_13_port, SUMB_12_12_port, SUMB_12_11_port, 
      SUMB_12_10_port, SUMB_12_9_port, SUMB_12_8_port, SUMB_12_7_port, 
      SUMB_12_6_port, SUMB_12_5_port, SUMB_12_4_port, SUMB_12_3_port, 
      SUMB_12_2_port, SUMB_12_1_port, SUMB_11_14_port, SUMB_11_13_port, 
      SUMB_11_12_port, SUMB_11_11_port, SUMB_11_10_port, SUMB_11_9_port, 
      SUMB_11_8_port, SUMB_11_7_port, SUMB_11_6_port, SUMB_11_5_port, 
      SUMB_11_4_port, SUMB_11_3_port, SUMB_11_2_port, SUMB_11_1_port, 
      SUMB_10_14_port, SUMB_10_13_port, SUMB_10_12_port, SUMB_10_11_port, 
      SUMB_10_10_port, SUMB_10_9_port, SUMB_10_8_port, SUMB_10_7_port, 
      SUMB_10_6_port, SUMB_10_5_port, SUMB_10_4_port, SUMB_10_3_port, 
      SUMB_10_2_port, SUMB_10_1_port, SUMB_9_14_port, SUMB_9_13_port, 
      SUMB_9_12_port, SUMB_9_11_port, SUMB_9_10_port, SUMB_9_9_port, 
      SUMB_9_8_port, SUMB_9_7_port, SUMB_9_6_port, SUMB_9_5_port, SUMB_9_4_port
      , SUMB_9_3_port, SUMB_9_2_port, SUMB_9_1_port, SUMB_8_14_port, 
      SUMB_8_13_port, SUMB_8_12_port, SUMB_8_11_port, SUMB_8_10_port, 
      SUMB_8_9_port, SUMB_8_8_port, SUMB_8_7_port, SUMB_8_6_port, SUMB_8_5_port
      , SUMB_8_4_port, SUMB_8_3_port, SUMB_8_2_port, SUMB_8_1_port, 
      SUMB_7_14_port, SUMB_7_13_port, SUMB_7_12_port, SUMB_7_11_port, 
      SUMB_7_10_port, SUMB_7_9_port, SUMB_7_8_port, SUMB_7_7_port, 
      SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, SUMB_7_3_port, SUMB_7_2_port
      , SUMB_7_1_port, SUMB_6_14_port, SUMB_6_13_port, SUMB_6_12_port, 
      SUMB_6_11_port, SUMB_6_10_port, SUMB_6_9_port, SUMB_6_8_port, 
      SUMB_6_7_port, SUMB_6_6_port, SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port
      , SUMB_6_2_port, SUMB_6_1_port, SUMB_5_14_port, SUMB_5_13_port, 
      SUMB_5_12_port, SUMB_5_11_port, SUMB_5_10_port, SUMB_5_9_port, 
      SUMB_5_8_port, SUMB_5_7_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port
      , SUMB_5_3_port, SUMB_5_2_port, SUMB_5_1_port, SUMB_4_14_port, 
      SUMB_4_13_port, SUMB_4_12_port, SUMB_4_11_port, SUMB_4_10_port, 
      SUMB_4_9_port, SUMB_4_8_port, SUMB_4_7_port, SUMB_4_6_port, SUMB_4_5_port
      , SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, 
      SUMB_3_14_port, SUMB_3_13_port, SUMB_3_12_port, SUMB_3_11_port, 
      SUMB_3_10_port, SUMB_3_9_port, SUMB_3_8_port, SUMB_3_7_port, 
      SUMB_3_6_port, SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port
      , SUMB_3_1_port, SUMB_2_14_port, SUMB_2_13_port, SUMB_2_12_port, 
      SUMB_2_11_port, SUMB_2_10_port, SUMB_2_9_port, SUMB_2_8_port, 
      SUMB_2_7_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, SUMB_1_14_port, SUMB_1_13_port, 
      SUMB_1_12_port, SUMB_1_11_port, SUMB_1_10_port, SUMB_1_9_port, 
      SUMB_1_8_port, SUMB_1_7_port, SUMB_1_6_port, SUMB_1_5_port, SUMB_1_4_port
      , SUMB_1_3_port, SUMB_1_2_port, SUMB_1_1_port, A1_28_port, A1_27_port, 
      A1_26_port, A1_25_port, A1_24_port, A1_23_port, A1_22_port, A1_21_port, 
      A1_20_port, A1_19_port, A1_18_port, A1_17_port, A1_16_port, A1_15_port, 
      A1_14_port, A1_13_port, A1_12_port, A1_11_port, A1_10_port, A1_9_port, 
      A1_8_port, A1_7_port, A1_6_port, A1_5_port, A1_4_port, A1_3_port, 
      A1_2_port, A1_1_port, A1_0_port, A2_21_port, A2_14_port, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, 
      n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, 
      n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_7 : FAX1 port map( A => ab_15_7_port, B => CARRYB_14_7_port, C => 
                           SUMB_14_8_port, YC => CARRYB_15_7_port, YS => 
                           SUMB_15_7_port);
   S4_8 : FAX1 port map( A => ab_15_8_port, B => CARRYB_14_8_port, C => 
                           SUMB_14_9_port, YC => CARRYB_15_8_port, YS => 
                           SUMB_15_8_port);
   S4_9 : FAX1 port map( A => ab_15_9_port, B => CARRYB_14_9_port, C => 
                           SUMB_14_10_port, YC => CARRYB_15_9_port, YS => 
                           SUMB_15_9_port);
   S4_10 : FAX1 port map( A => ab_15_10_port, B => CARRYB_14_10_port, C => 
                           SUMB_14_11_port, YC => CARRYB_15_10_port, YS => 
                           SUMB_15_10_port);
   S4_11 : FAX1 port map( A => ab_15_11_port, B => CARRYB_14_11_port, C => 
                           SUMB_14_12_port, YC => CARRYB_15_11_port, YS => 
                           SUMB_15_11_port);
   S4_12 : FAX1 port map( A => ab_15_12_port, B => CARRYB_14_12_port, C => 
                           SUMB_14_13_port, YC => CARRYB_15_12_port, YS => 
                           SUMB_15_12_port);
   S4_13 : FAX1 port map( A => ab_15_13_port, B => CARRYB_14_13_port, C => 
                           SUMB_14_14_port, YC => CARRYB_15_13_port, YS => 
                           SUMB_15_13_port);
   S5_14 : FAX1 port map( A => ab_15_14_port, B => CARRYB_14_14_port, C => 
                           ab_14_15_port, YC => CARRYB_15_14_port, YS => 
                           SUMB_15_14_port);
   S14_15 : FAX1 port map( A => n1096, B => n1095, C => ab_15_15_port, YC => 
                           CARRYB_15_15_port, YS => SUMB_15_15_port);
   S2_14_9 : FAX1 port map( A => ab_14_9_port, B => CARRYB_13_9_port, C => 
                           SUMB_13_10_port, YC => CARRYB_14_9_port, YS => 
                           SUMB_14_9_port);
   S2_14_10 : FAX1 port map( A => ab_14_10_port, B => CARRYB_13_10_port, C => 
                           SUMB_13_11_port, YC => CARRYB_14_10_port, YS => 
                           SUMB_14_10_port);
   S2_14_11 : FAX1 port map( A => ab_14_11_port, B => CARRYB_13_11_port, C => 
                           SUMB_13_12_port, YC => CARRYB_14_11_port, YS => 
                           SUMB_14_11_port);
   S2_14_12 : FAX1 port map( A => ab_14_12_port, B => CARRYB_13_12_port, C => 
                           SUMB_13_13_port, YC => CARRYB_14_12_port, YS => 
                           SUMB_14_12_port);
   S2_14_13 : FAX1 port map( A => ab_14_13_port, B => CARRYB_13_13_port, C => 
                           SUMB_13_14_port, YC => CARRYB_14_13_port, YS => 
                           SUMB_14_13_port);
   S3_14_14 : FAX1 port map( A => ab_14_14_port, B => CARRYB_13_14_port, C => 
                           ab_13_15_port, YC => CARRYB_14_14_port, YS => 
                           SUMB_14_14_port);
   S2_13_10 : FAX1 port map( A => ab_13_10_port, B => CARRYB_12_10_port, C => 
                           SUMB_12_11_port, YC => CARRYB_13_10_port, YS => 
                           SUMB_13_10_port);
   S2_13_11 : FAX1 port map( A => ab_13_11_port, B => CARRYB_12_11_port, C => 
                           SUMB_12_12_port, YC => CARRYB_13_11_port, YS => 
                           SUMB_13_11_port);
   S2_13_12 : FAX1 port map( A => ab_13_12_port, B => CARRYB_12_12_port, C => 
                           SUMB_12_13_port, YC => CARRYB_13_12_port, YS => 
                           SUMB_13_12_port);
   S2_13_13 : FAX1 port map( A => ab_13_13_port, B => CARRYB_12_13_port, C => 
                           SUMB_12_14_port, YC => CARRYB_13_13_port, YS => 
                           SUMB_13_13_port);
   S3_13_14 : FAX1 port map( A => ab_13_14_port, B => CARRYB_12_14_port, C => 
                           ab_12_15_port, YC => CARRYB_13_14_port, YS => 
                           SUMB_13_14_port);
   S2_12_8 : FAX1 port map( A => ab_12_8_port, B => CARRYB_11_8_port, C => 
                           SUMB_11_9_port, YC => CARRYB_12_8_port, YS => 
                           SUMB_12_8_port);
   S2_12_10 : FAX1 port map( A => ab_12_10_port, B => CARRYB_11_10_port, C => 
                           SUMB_11_11_port, YC => CARRYB_12_10_port, YS => 
                           SUMB_12_10_port);
   S2_12_11 : FAX1 port map( A => ab_12_11_port, B => CARRYB_11_11_port, C => 
                           SUMB_11_12_port, YC => CARRYB_12_11_port, YS => 
                           SUMB_12_11_port);
   S2_12_12 : FAX1 port map( A => ab_12_12_port, B => CARRYB_11_12_port, C => 
                           SUMB_11_13_port, YC => CARRYB_12_12_port, YS => 
                           SUMB_12_12_port);
   S2_12_13 : FAX1 port map( A => ab_12_13_port, B => CARRYB_11_13_port, C => 
                           SUMB_11_14_port, YC => CARRYB_12_13_port, YS => 
                           SUMB_12_13_port);
   S3_12_14 : FAX1 port map( A => ab_12_14_port, B => CARRYB_11_14_port, C => 
                           ab_11_15_port, YC => CARRYB_12_14_port, YS => 
                           SUMB_12_14_port);
   S2_11_11 : FAX1 port map( A => ab_11_11_port, B => CARRYB_10_11_port, C => 
                           SUMB_10_12_port, YC => CARRYB_11_11_port, YS => 
                           SUMB_11_11_port);
   S2_11_12 : FAX1 port map( A => ab_11_12_port, B => CARRYB_10_12_port, C => 
                           SUMB_10_13_port, YC => CARRYB_11_12_port, YS => 
                           SUMB_11_12_port);
   S2_11_13 : FAX1 port map( A => ab_11_13_port, B => CARRYB_10_13_port, C => 
                           SUMB_10_14_port, YC => CARRYB_11_13_port, YS => 
                           SUMB_11_13_port);
   S3_11_14 : FAX1 port map( A => ab_11_14_port, B => CARRYB_10_14_port, C => 
                           ab_10_15_port, YC => CARRYB_11_14_port, YS => 
                           SUMB_11_14_port);
   S1_10_0 : FAX1 port map( A => ab_10_0_port, B => SUMB_9_1_port, C => 
                           CARRYB_9_0_port, YC => CARRYB_10_0_port, YS => 
                           A1_8_port);
   S2_10_13 : FAX1 port map( A => ab_10_13_port, B => CARRYB_9_13_port, C => 
                           SUMB_9_14_port, YC => CARRYB_10_13_port, YS => 
                           SUMB_10_13_port);
   S3_10_14 : FAX1 port map( A => ab_10_14_port, B => CARRYB_9_14_port, C => 
                           ab_9_15_port, YC => CARRYB_10_14_port, YS => 
                           SUMB_10_14_port);
   S2_9_1 : FAX1 port map( A => ab_9_1_port, B => CARRYB_8_1_port, C => 
                           SUMB_8_2_port, YC => CARRYB_9_1_port, YS => 
                           SUMB_9_1_port);
   S2_9_11 : FAX1 port map( A => CARRYB_8_11_port, B => ab_9_11_port, C => 
                           SUMB_8_12_port, YC => CARRYB_9_11_port, YS => 
                           SUMB_9_11_port);
   S3_9_14 : FAX1 port map( A => ab_9_14_port, B => CARRYB_8_14_port, C => 
                           ab_8_15_port, YC => CARRYB_9_14_port, YS => 
                           SUMB_9_14_port);
   S2_8_12 : FAX1 port map( A => ab_8_12_port, B => CARRYB_7_12_port, C => 
                           SUMB_7_13_port, YC => CARRYB_8_12_port, YS => 
                           SUMB_8_12_port);
   S2_8_13 : FAX1 port map( A => ab_8_13_port, B => CARRYB_7_13_port, C => 
                           SUMB_7_14_port, YC => CARRYB_8_13_port, YS => 
                           SUMB_8_13_port);
   S3_8_14 : FAX1 port map( A => ab_8_14_port, B => CARRYB_7_14_port, C => 
                           ab_7_15_port, YC => CARRYB_8_14_port, YS => 
                           SUMB_8_14_port);
   S2_7_11 : FAX1 port map( A => ab_7_11_port, B => n251, C => SUMB_6_12_port, 
                           YC => CARRYB_7_11_port, YS => SUMB_7_11_port);
   S3_7_14 : FAX1 port map( A => ab_7_14_port, B => CARRYB_6_14_port, C => 
                           ab_6_15_port, YC => CARRYB_7_14_port, YS => 
                           SUMB_7_14_port);
   S1_6_0 : FAX1 port map( A => CARRYB_5_0_port, B => ab_6_0_port, C => 
                           SUMB_5_1_port, YC => CARRYB_6_0_port, YS => 
                           A1_4_port);
   S1_5_0 : FAX1 port map( A => CARRYB_4_0_port, B => ab_5_0_port, C => 
                           SUMB_4_1_port, YC => CARRYB_5_0_port, YS => 
                           A1_3_port);
   S3_5_14 : FAX1 port map( A => ab_5_14_port, B => CARRYB_4_14_port, C => 
                           ab_4_15_port, YC => CARRYB_5_14_port, YS => 
                           SUMB_5_14_port);
   S1_4_0 : FAX1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, C => 
                           SUMB_3_1_port, YC => CARRYB_4_0_port, YS => 
                           A1_2_port);
   S3_3_14 : FAX1 port map( A => ab_3_14_port, B => ab_2_15_port, C => 
                           CARRYB_2_14_port, YC => CARRYB_3_14_port, YS => 
                           SUMB_3_14_port);
   S1_2_0 : FAX1 port map( A => ab_2_0_port, B => n1020, C => SUMB_1_1_port, YC
                           => CARRYB_2_0_port, YS => A1_0_port);
   FS_1 : matrix_math_DW01_add_23 port map( A(29) => n1094, A(28) => A1_28_port
                           , A(27) => A1_27_port, A(26) => A1_26_port, A(25) =>
                           A1_25_port, A(24) => A1_24_port, A(23) => A1_23_port
                           , A(22) => A1_22_port, A(21) => A1_21_port, A(20) =>
                           A1_20_port, A(19) => A1_19_port, A(18) => A1_18_port
                           , A(17) => A1_17_port, A(16) => A1_16_port, A(15) =>
                           A1_15_port, A(14) => A1_14_port, A(13) => A1_13_port
                           , A(12) => A1_12_port, A(11) => A1_11_port, A(10) =>
                           A1_10_port, A(9) => A1_9_port, A(8) => A1_8_port, 
                           A(7) => A1_7_port, A(6) => A1_6_port, A(5) => 
                           A1_5_port, A(4) => A1_4_port, A(3) => A1_3_port, 
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(29) => n95, B(28) => n94, B(27) => n93,
                           B(26) => n92, B(25) => n91, B(24) => n90, B(23) => 
                           n89, B(22) => n88, B(21) => A2_21_port, B(20) => 
                           n1019, B(19) => n1018, B(18) => n1017, B(17) => 
                           n1016, B(16) => n1015, B(15) => n1014, B(14) => 
                           A2_14_port, B(13) => n1099, B(12) => n1099, B(11) =>
                           n1099, B(10) => n1099, B(9) => n1099, B(8) => n1099,
                           B(7) => n1099, B(6) => n1099, B(5) => n1099, B(4) =>
                           n1099, B(3) => n1099, B(2) => n1099, B(1) => n1099, 
                           B(0) => X_Logic0_port, CI => X_Logic0_port, SUM(29) 
                           => n_1177, SUM(28) => n_1178, SUM(27) => n_1179, 
                           SUM(26) => n_1180, SUM(25) => n_1181, SUM(24) => 
                           n_1182, SUM(23) => n_1183, SUM(22) => n_1184, 
                           SUM(21) => PRODUCT(23), SUM(20) => PRODUCT(22), 
                           SUM(19) => PRODUCT(21), SUM(18) => PRODUCT(20), 
                           SUM(17) => PRODUCT(19), SUM(16) => PRODUCT(18), 
                           SUM(15) => PRODUCT(17), SUM(14) => PRODUCT(16), 
                           SUM(13) => PRODUCT(15), SUM(12) => PRODUCT(14), 
                           SUM(11) => PRODUCT(13), SUM(10) => PRODUCT(12), 
                           SUM(9) => PRODUCT(11), SUM(8) => PRODUCT(10), SUM(7)
                           => PRODUCT(9), SUM(6) => PRODUCT(8), SUM(5) => 
                           PRODUCT(7), SUM(4) => PRODUCT(6), SUM(3) => 
                           PRODUCT(5), SUM(2) => PRODUCT(4), SUM(1) => 
                           PRODUCT(3), SUM(0) => PRODUCT(2), CO => n_1185);
   U2 : AND2X2 port map( A => ab_1_8_port, B => ab_0_9_port, Y => n3);
   U3 : BUFX2 port map( A => n739, Y => n4);
   U4 : NAND3X1 port map( A => n670, B => n669, C => n668, Y => n5);
   U5 : BUFX2 port map( A => n741, Y => n6);
   U6 : NAND3X1 port map( A => n820, B => n821, C => n822, Y => n7);
   U7 : BUFX2 port map( A => n603, Y => n8);
   U8 : XOR2X1 port map( A => n62, B => n9, Y => SUMB_3_11_port);
   U9 : XNOR2X1 port map( A => CARRYB_2_11_port, B => ab_3_11_port, Y => n9);
   U10 : XNOR2X1 port map( A => n10, B => n11, Y => SUMB_6_4_port);
   U11 : XOR2X1 port map( A => SUMB_5_5_port, B => ab_6_4_port, Y => n10);
   U12 : INVX1 port map( A => CARRYB_5_4_port, Y => n11);
   U13 : BUFX2 port map( A => n187, Y => n12);
   U14 : XOR2X1 port map( A => n13, B => n36, Y => SUMB_13_1_port);
   U15 : XOR2X1 port map( A => CARRYB_12_1_port, B => n271, Y => n13);
   U16 : INVX1 port map( A => SUMB_12_2_port, Y => n36);
   U17 : INVX2 port map( A => n913, Y => n914);
   U18 : XOR2X1 port map( A => n14, B => ab_2_9_port, Y => n15);
   U19 : NAND2X1 port map( A => ab_0_10_port, B => n429, Y => n14);
   U20 : XNOR2X1 port map( A => n15, B => SUMB_1_10_port, Y => SUMB_2_9_port);
   U21 : BUFX2 port map( A => n896, Y => n16);
   U22 : BUFX2 port map( A => SUMB_5_2_port, Y => n17);
   U23 : XOR2X1 port map( A => CARRYB_9_5_port, B => ab_10_5_port, Y => n281);
   U24 : NAND2X1 port map( A => ab_8_3_port, B => n141, Y => n18);
   U25 : XOR2X1 port map( A => CARRYB_11_4_port, B => ab_12_4_port, Y => n47);
   U26 : BUFX2 port map( A => SUMB_10_11_port, Y => n19);
   U27 : BUFX2 port map( A => n188, Y => n20);
   U28 : XNOR2X1 port map( A => n21, B => n218, Y => SUMB_5_8_port);
   U29 : XOR2X1 port map( A => CARRYB_4_8_port, B => ab_5_8_port, Y => n21);
   U30 : XNOR2X1 port map( A => n22, B => n45, Y => SUMB_7_7_port);
   U31 : XOR2X1 port map( A => CARRYB_6_7_port, B => ab_7_7_port, Y => n22);
   U32 : XNOR2X1 port map( A => CARRYB_2_9_port, B => n23, Y => n182);
   U33 : INVX8 port map( A => ab_3_9_port, Y => n23);
   U34 : BUFX2 port map( A => n958, Y => n24);
   U35 : INVX2 port map( A => SUMB_4_5_port, Y => n527);
   U36 : INVX2 port map( A => SUMB_6_3_port, Y => n453);
   U37 : XNOR2X1 port map( A => n25, B => SUMB_9_7_port, Y => SUMB_10_6_port);
   U38 : XNOR2X1 port map( A => CARRYB_9_6_port, B => ab_10_6_port, Y => n25);
   U39 : XNOR2X1 port map( A => n26, B => SUMB_6_9_port, Y => SUMB_7_8_port);
   U40 : XNOR2X1 port map( A => CARRYB_6_8_port, B => n40, Y => n26);
   U41 : BUFX2 port map( A => n787, Y => n27);
   U42 : XNOR2X1 port map( A => n235, B => n179, Y => n28);
   U43 : XNOR2X1 port map( A => n29, B => SUMB_9_5_port, Y => SUMB_10_4_port);
   U44 : XNOR2X1 port map( A => CARRYB_9_4_port, B => ab_10_4_port, Y => n29);
   U45 : XNOR2X1 port map( A => n30, B => SUMB_13_6_port, Y => SUMB_14_5_port);
   U46 : XNOR2X1 port map( A => CARRYB_13_5_port, B => n48, Y => n30);
   U47 : XOR2X1 port map( A => n454, B => n31, Y => n227);
   U48 : INVX8 port map( A => ab_12_3_port, Y => n31);
   U49 : BUFX2 port map( A => SUMB_12_1_port, Y => n32);
   U50 : XOR2X1 port map( A => n394, B => n33, Y => n432);
   U51 : INVX8 port map( A => ab_14_2_port, Y => n33);
   U52 : XOR2X1 port map( A => CARRYB_8_3_port, B => n34, Y => n724);
   U53 : INVX8 port map( A => ab_9_3_port, Y => n34);
   U54 : XOR2X1 port map( A => n35, B => n76, Y => SUMB_9_5_port);
   U55 : XOR2X1 port map( A => CARRYB_8_5_port, B => ab_9_5_port, Y => n35);
   U56 : XOR2X1 port map( A => CARRYB_11_5_port, B => n37, Y => n132);
   U57 : INVX8 port map( A => ab_12_5_port, Y => n37);
   U58 : XOR2X1 port map( A => n38, B => SUMB_4_8_port, Y => SUMB_5_7_port);
   U59 : XOR2X1 port map( A => CARRYB_4_7_port, B => ab_5_7_port, Y => n38);
   U60 : BUFX2 port map( A => n959, Y => n39);
   U61 : INVX8 port map( A => n526, Y => n40);
   U62 : XNOR2X1 port map( A => n41, B => SUMB_5_9_port, Y => SUMB_6_8_port);
   U63 : XNOR2X1 port map( A => CARRYB_5_8_port, B => ab_6_8_port, Y => n41);
   U64 : BUFX2 port map( A => A(1), Y => n42);
   U65 : INVX1 port map( A => A(1), Y => n430);
   U66 : BUFX2 port map( A => SUMB_2_14_port, Y => n43);
   U67 : BUFX2 port map( A => SUMB_4_13_port, Y => n44);
   U68 : INVX2 port map( A => SUMB_4_9_port, Y => n218);
   U69 : INVX2 port map( A => SUMB_6_8_port, Y => n45);
   U70 : XOR2X1 port map( A => n46, B => CARRYB_11_6_port, Y => SUMB_12_6_port)
                           ;
   U71 : XNOR2X1 port map( A => SUMB_11_7_port, B => n355, Y => n46);
   U72 : XOR2X1 port map( A => n47, B => SUMB_11_5_port, Y => SUMB_12_4_port);
   U73 : INVX8 port map( A => n397, Y => n48);
   U74 : XOR2X1 port map( A => n49, B => n511, Y => SUMB_2_14_port);
   U75 : XNOR2X1 port map( A => n196, B => ab_2_14_port, Y => n49);
   U76 : INVX4 port map( A => B(13), Y => n1057);
   U77 : XNOR2X1 port map( A => n50, B => SUMB_1_13_port, Y => SUMB_2_12_port);
   U78 : XNOR2X1 port map( A => n388, B => ab_2_12_port, Y => n50);
   U79 : XNOR2X1 port map( A => CARRYB_14_3_port, B => n80, Y => n146);
   U80 : BUFX2 port map( A => n872, Y => n51);
   U81 : XNOR2X1 port map( A => n835, B => n52, Y => n541);
   U82 : INVX8 port map( A => ab_6_9_port, Y => n52);
   U83 : XNOR2X1 port map( A => n53, B => SUMB_10_8_port, Y => SUMB_11_7_port);
   U84 : XOR2X1 port map( A => CARRYB_10_7_port, B => n654, Y => n53);
   U85 : XNOR2X1 port map( A => n54, B => SUMB_14_6_port, Y => SUMB_15_5_port);
   U86 : XNOR2X1 port map( A => CARRYB_14_5_port, B => ab_15_5_port, Y => n54);
   U87 : XOR2X1 port map( A => n182, B => n68, Y => n55);
   U88 : NAND3X1 port map( A => n598, B => n599, C => n600, Y => n56);
   U89 : INVX2 port map( A => SUMB_12_4_port, Y => n387);
   U90 : BUFX2 port map( A => n899, Y => n57);
   U91 : XNOR2X1 port map( A => CARRYB_7_6_port, B => n58, Y => n107);
   U92 : INVX8 port map( A => n224, Y => n58);
   U93 : INVX2 port map( A => SUMB_2_11_port, Y => n59);
   U94 : INVX2 port map( A => n59, Y => n60);
   U95 : XOR2X1 port map( A => n61, B => SUMB_1_12_port, Y => SUMB_2_11_port);
   U96 : XNOR2X1 port map( A => n174, B => ab_2_11_port, Y => n61);
   U97 : INVX1 port map( A => SUMB_2_12_port, Y => n62);
   U98 : XNOR2X1 port map( A => CARRYB_13_3_port, B => n474, Y => n63);
   U99 : XOR2X1 port map( A => n797, B => n64, Y => n386);
   U100 : INVX8 port map( A => n73, Y => n64);
   U101 : XOR2X1 port map( A => n65, B => SUMB_4_10_port, Y => SUMB_5_9_port);
   U102 : XNOR2X1 port map( A => CARRYB_4_9_port, B => n173, Y => n65);
   U103 : INVX4 port map( A => B(15), Y => n1095);
   U104 : XNOR2X1 port map( A => n66, B => SUMB_5_13_port, Y => SUMB_6_12_port)
                           ;
   U105 : XNOR2X1 port map( A => ab_6_12_port, B => CARRYB_5_12_port, Y => n66)
                           ;
   U106 : AND2X1 port map( A => SUMB_15_6_port, B => CARRYB_15_5_port, Y => 
                           n1019);
   U107 : XOR2X1 port map( A => n67, B => n276, Y => SUMB_12_1_port);
   U108 : XOR2X1 port map( A => n666, B => ab_12_1_port, Y => n67);
   U109 : XOR2X1 port map( A => n216, B => n272, Y => n68);
   U110 : AND2X2 port map( A => ab_0_10_port, B => n429, Y => n69);
   U111 : XOR2X1 port map( A => CARRYB_10_4_port, B => n70, Y => n240);
   U112 : INVX8 port map( A => ab_11_4_port, Y => n70);
   U113 : XOR2X1 port map( A => CARRYB_14_2_port, B => n71, Y => n255);
   U114 : INVX8 port map( A => n72, Y => n71);
   U115 : INVX8 port map( A => ab_15_2_port, Y => n72);
   U116 : INVX8 port map( A => ab_13_3_port, Y => n73);
   U117 : BUFX2 port map( A => SUMB_9_4_port, Y => n74);
   U118 : XOR2X1 port map( A => CARRYB_12_2_port, B => n75, Y => n164);
   U119 : INVX8 port map( A => ab_13_2_port, Y => n75);
   U120 : XOR2X1 port map( A => n107, B => n217, Y => n76);
   U121 : XOR2X1 port map( A => n123, B => n121, Y => n77);
   U122 : INVX4 port map( A => n1053, Y => n1054);
   U123 : INVX1 port map( A => B(11), Y => n1053);
   U124 : AND2X2 port map( A => ab_0_3_port, B => n1022, Y => n78);
   U125 : AND2X2 port map( A => ab_0_4_port, B => ab_1_3_port, Y => n1021);
   U126 : XOR2X1 port map( A => SUMB_7_9_port, B => n79, Y => n81);
   U127 : INVX8 port map( A => n211, Y => n79);
   U128 : INVX8 port map( A => ab_15_3_port, Y => n80);
   U129 : XOR2X1 port map( A => n81, B => CARRYB_7_8_port, Y => SUMB_8_8_port);
   U130 : XOR2X1 port map( A => n181, B => n356, Y => n82);
   U131 : XOR2X1 port map( A => SUMB_5_12_port, B => ab_6_11_port, Y => n83);
   U132 : XOR2X1 port map( A => n83, B => CARRYB_5_11_port, Y => SUMB_6_11_port
                           );
   U133 : NAND2X1 port map( A => CARRYB_5_11_port, B => SUMB_5_12_port, Y => 
                           n84);
   U134 : NAND2X1 port map( A => CARRYB_5_11_port, B => ab_6_11_port, Y => n85)
                           ;
   U135 : NAND2X1 port map( A => SUMB_5_12_port, B => ab_6_11_port, Y => n86);
   U136 : NAND3X1 port map( A => n85, B => n84, C => n86, Y => CARRYB_6_11_port
                           );
   U137 : INVX2 port map( A => SUMB_7_6_port, Y => n235);
   U138 : XOR2X1 port map( A => CARRYB_5_7_port, B => n87, Y => n715);
   U139 : INVX8 port map( A => ab_6_7_port, Y => n87);
   U140 : INVX2 port map( A => ab_10_7_port, Y => n119);
   U141 : INVX2 port map( A => ab_10_3_port, Y => n577);
   U142 : INVX2 port map( A => ab_5_9_port, Y => n173);
   U143 : INVX2 port map( A => ab_5_10_port, Y => n213);
   U144 : INVX2 port map( A => ab_5_6_port, Y => n532);
   U145 : INVX2 port map( A => ab_4_6_port, Y => n208);
   U146 : INVX2 port map( A => ab_8_8_port, Y => n211);
   U147 : INVX2 port map( A => ab_13_3_port, Y => n520);
   U148 : INVX2 port map( A => ab_12_6_port, Y => n355);
   U149 : INVX2 port map( A => ab_10_2_port, Y => n731);
   U150 : INVX2 port map( A => ab_12_2_port, Y => n448);
   U151 : INVX2 port map( A => ab_7_8_port, Y => n526);
   U152 : INVX2 port map( A => ab_7_9_port, Y => n234);
   U153 : INVX2 port map( A => ab_6_6_port, Y => n228);
   U154 : INVX2 port map( A => ab_6_5_port, Y => n150);
   U155 : INVX2 port map( A => ab_5_5_port, Y => n434);
   U156 : INVX2 port map( A => ab_8_6_port, Y => n224);
   U157 : INVX2 port map( A => ab_14_3_port, Y => n474);
   U158 : INVX2 port map( A => ab_13_4_port, Y => n590);
   U159 : INVX2 port map( A => ab_8_2_port, Y => n463);
   U160 : INVX2 port map( A => n1034, Y => n1035);
   U161 : INVX2 port map( A => ab_14_5_port, Y => n397);
   U162 : INVX2 port map( A => ab_15_6_port, Y => n540);
   U163 : INVX2 port map( A => n1080, Y => n1081);
   U164 : INVX2 port map( A => ab_13_1_port, Y => n271);
   U165 : INVX2 port map( A => ab_11_10_port, Y => n197);
   U166 : INVX2 port map( A => n1046, Y => n1047);
   U167 : AND2X2 port map( A => SUMB_15_8_port, B => CARRYB_15_7_port, Y => n88
                           );
   U168 : AND2X2 port map( A => SUMB_15_9_port, B => CARRYB_15_8_port, Y => n89
                           );
   U169 : AND2X2 port map( A => SUMB_15_10_port, B => CARRYB_15_9_port, Y => 
                           n90);
   U170 : AND2X2 port map( A => SUMB_15_11_port, B => CARRYB_15_10_port, Y => 
                           n91);
   U171 : AND2X2 port map( A => SUMB_15_12_port, B => CARRYB_15_11_port, Y => 
                           n92);
   U172 : AND2X2 port map( A => SUMB_15_13_port, B => CARRYB_15_12_port, Y => 
                           n93);
   U173 : AND2X2 port map( A => SUMB_15_14_port, B => CARRYB_15_13_port, Y => 
                           n94);
   U174 : AND2X2 port map( A => SUMB_15_15_port, B => CARRYB_15_14_port, Y => 
                           n95);
   U175 : AND2X2 port map( A => ab_0_2_port, B => ab_1_1_port, Y => n96);
   U176 : AND2X2 port map( A => ab_0_5_port, B => ab_1_4_port, Y => n97);
   U177 : INVX2 port map( A => n169, Y => n104);
   U178 : AND2X1 port map( A => n789, B => n791, Y => n98);
   U179 : AND2X1 port map( A => n381, B => n380, Y => n99);
   U180 : INVX2 port map( A => ab_11_3_port, Y => n464);
   U181 : BUFX2 port map( A => SUMB_4_7_port, Y => n100);
   U182 : BUFX2 port map( A => SUMB_5_6_port, Y => n101);
   U183 : XOR2X1 port map( A => SUMB_3_11_port, B => n102, Y => SUMB_4_10_port)
                           ;
   U184 : XOR2X1 port map( A => CARRYB_3_10_port, B => ab_4_10_port, Y => n102)
                           ;
   U185 : INVX2 port map( A => n1061, Y => n103);
   U186 : INVX4 port map( A => n1061, Y => n1062);
   U187 : INVX1 port map( A => SUMB_11_2_port, Y => n276);
   U188 : INVX2 port map( A => ab_2_10_port, Y => n169);
   U189 : INVX1 port map( A => n1061, Y => n105);
   U190 : BUFX2 port map( A => ab_2_11_port, Y => n106);
   U191 : XOR2X1 port map( A => n107, B => n217, Y => SUMB_8_6_port);
   U192 : INVX1 port map( A => SUMB_10_3_port, Y => n149);
   U193 : AND2X2 port map( A => n42, B => n1045, Y => ab_1_6_port);
   U194 : AND2X1 port map( A => n983, B => B(1), Y => ab_1_1_port);
   U195 : NAND3X1 port map( A => n368, B => n367, C => n369, Y => n108);
   U196 : NAND3X1 port map( A => n881, B => n882, C => n883, Y => n109);
   U197 : BUFX2 port map( A => n845, Y => n110);
   U198 : NAND3X1 port map( A => n496, B => n497, C => n498, Y => n111);
   U199 : XNOR2X1 port map( A => n112, B => SUMB_10_4_port, Y => SUMB_11_3_port
                           );
   U200 : XNOR2X1 port map( A => n1028, B => n464, Y => n112);
   U201 : AND2X1 port map( A => ab_1_11_port, B => ab_0_12_port, Y => n186);
   U202 : BUFX2 port map( A => SUMB_15_0_port, Y => n113);
   U203 : INVX1 port map( A => CARRYB_15_0_port, Y => n114);
   U204 : INVX1 port map( A => n114, Y => n115);
   U205 : NAND3X1 port map( A => n12, B => n20, C => n189, Y => n116);
   U206 : BUFX2 port map( A => n873, Y => n117);
   U207 : XOR2X1 port map( A => n118, B => SUMB_5_7_port, Y => SUMB_6_6_port);
   U208 : XNOR2X1 port map( A => CARRYB_5_6_port, B => n228, Y => n118);
   U209 : XOR2X1 port map( A => CARRYB_9_7_port, B => n119, Y => n273);
   U210 : XOR2X1 port map( A => n255, B => n183, Y => SUMB_15_2_port);
   U211 : NAND3X1 port map( A => n385, B => n384, C => n383, Y => 
                           CARRYB_2_11_port);
   U212 : XNOR2X1 port map( A => n1025, B => ab_2_13_port, Y => n779);
   U213 : NAND3X1 port map( A => n554, B => n556, C => n555, Y => n394);
   U214 : BUFX2 port map( A => n846, Y => n120);
   U215 : XNOR2X1 port map( A => n164, B => n200, Y => n121);
   U216 : XOR2X1 port map( A => n589, B => n122, Y => SUMB_8_4_port);
   U217 : XNOR2X1 port map( A => CARRYB_7_4_port, B => ab_8_4_port, Y => n122);
   U218 : XOR2X1 port map( A => n123, B => n121, Y => SUMB_14_1_port);
   U219 : XNOR2X1 port map( A => n1030, B => ab_14_1_port, Y => n123);
   U220 : NAND3X1 port map( A => n716, B => n717, C => n718, Y => n124);
   U221 : NAND3X1 port map( A => n844, B => n110, C => n120, Y => n125);
   U222 : XOR2X1 port map( A => n724, B => n329, Y => n126);
   U223 : XNOR2X1 port map( A => n127, B => n28, Y => SUMB_9_4_port);
   U224 : XNOR2X1 port map( A => CARRYB_8_4_port, B => ab_9_4_port, Y => n127);
   U225 : NAND3X1 port map( A => n823, B => n824, C => n825, Y => n128);
   U226 : NAND3X1 port map( A => n891, B => n892, C => n893, Y => n129);
   U227 : NAND3X1 port map( A => n338, B => n337, C => n339, Y => n130);
   U228 : BUFX2 port map( A => n751, Y => n131);
   U229 : XNOR2X1 port map( A => n132, B => SUMB_11_6_port, Y => SUMB_12_5_port
                           );
   U230 : XNOR2X1 port map( A => n133, B => SUMB_10_7_port, Y => SUMB_11_6_port
                           );
   U231 : XNOR2X1 port map( A => CARRYB_10_6_port, B => ab_11_6_port, Y => n133
                           );
   U232 : NAND3X1 port map( A => n535, B => n533, C => n534, Y => n134);
   U233 : NAND3X1 port map( A => n331, B => n332, C => n333, Y => n135);
   U234 : NAND3X1 port map( A => n743, B => n744, C => n745, Y => n136);
   U235 : XOR2X1 port map( A => n432, B => n433, Y => n137);
   U236 : NAND3X1 port map( A => n515, B => n516, C => n517, Y => n138);
   U237 : BUFX2 port map( A => CARRYB_15_2_port, Y => n139);
   U238 : NAND3X1 port map( A => n606, B => n605, C => n607, Y => n140);
   U239 : NAND3X1 port map( A => n725, B => n727, C => n726, Y => n141);
   U240 : NAND3X1 port map( A => n598, B => n599, C => n600, Y => n142);
   U241 : NAND3X1 port map( A => n904, B => n906, C => n905, Y => n143);
   U242 : NAND3X1 port map( A => n635, B => n637, C => n636, Y => n144);
   U243 : NAND3X1 port map( A => n989, B => n990, C => n991, Y => n145);
   U244 : XOR2X1 port map( A => n146, B => SUMB_14_4_port, Y => SUMB_15_3_port)
                           ;
   U245 : XOR2X1 port map( A => n147, B => n575, Y => SUMB_7_4_port);
   U246 : XOR2X1 port map( A => CARRYB_6_4_port, B => ab_7_4_port, Y => n147);
   U247 : XOR2X1 port map( A => n545, B => ab_11_2_port, Y => n148);
   U248 : XNOR2X1 port map( A => n148, B => n149, Y => SUMB_11_2_port);
   U249 : XOR2X1 port map( A => CARRYB_5_5_port, B => n150, Y => n167);
   U250 : XOR2X1 port map( A => CARRYB_14_1_port, B => ab_15_1_port, Y => n547)
                           ;
   U251 : XNOR2X1 port map( A => n151, B => SUMB_8_8_port, Y => SUMB_9_7_port);
   U252 : XNOR2X1 port map( A => CARRYB_8_7_port, B => ab_9_7_port, Y => n151);
   U253 : XOR2X1 port map( A => n152, B => SUMB_6_6_port, Y => SUMB_7_5_port);
   U254 : XOR2X1 port map( A => CARRYB_6_5_port, B => ab_7_5_port, Y => n152);
   U255 : BUFX2 port map( A => n1065, Y => n153);
   U256 : XOR2X1 port map( A => ab_13_9_port, B => CARRYB_12_9_port, Y => n154)
                           ;
   U257 : XOR2X1 port map( A => n154, B => SUMB_12_10_port, Y => SUMB_13_9_port
                           );
   U258 : XOR2X1 port map( A => ab_14_8_port, B => CARRYB_13_8_port, Y => n155)
                           ;
   U259 : XOR2X1 port map( A => n155, B => SUMB_13_9_port, Y => SUMB_14_8_port)
                           ;
   U260 : NAND2X1 port map( A => ab_13_9_port, B => CARRYB_12_9_port, Y => n156
                           );
   U261 : NAND2X1 port map( A => ab_13_9_port, B => SUMB_12_10_port, Y => n157)
                           ;
   U262 : NAND2X1 port map( A => CARRYB_12_9_port, B => SUMB_12_10_port, Y => 
                           n158);
   U263 : NAND3X1 port map( A => n156, B => n157, C => n158, Y => 
                           CARRYB_13_9_port);
   U264 : NAND2X1 port map( A => ab_14_8_port, B => n108, Y => n159);
   U265 : NAND2X1 port map( A => ab_14_8_port, B => SUMB_13_9_port, Y => n160);
   U266 : NAND2X1 port map( A => n108, B => SUMB_13_9_port, Y => n161);
   U267 : NAND3X1 port map( A => n159, B => n160, C => n161, Y => 
                           CARRYB_14_8_port);
   U268 : BUFX2 port map( A => SUMB_3_13_port, Y => n162);
   U269 : NAND3X1 port map( A => n782, B => n780, C => n781, Y => n163);
   U270 : XNOR2X1 port map( A => n164, B => n200, Y => SUMB_13_2_port);
   U271 : BUFX2 port map( A => CARRYB_4_7_port, Y => n165);
   U272 : XNOR2X1 port map( A => n166, B => ab_1_8_port, Y => SUMB_1_8_port);
   U273 : NAND2X1 port map( A => B(9), B => n1062, Y => n166);
   U274 : XNOR2X1 port map( A => n167, B => n101, Y => SUMB_6_5_port);
   U275 : INVX1 port map( A => SUMB_3_7_port, Y => n254);
   U276 : XNOR2X1 port map( A => n168, B => n314, Y => SUMB_4_9_port);
   U277 : XOR2X1 port map( A => CARRYB_3_9_port, B => ab_4_9_port, Y => n168);
   U278 : BUFX2 port map( A => n466, Y => n170);
   U279 : XNOR2X1 port map( A => CARRYB_9_8_port, B => ab_10_8_port, Y => n357)
                           ;
   U280 : INVX2 port map( A => SUMB_2_13_port, Y => n356);
   U281 : INVX2 port map( A => CARRYB_3_7_port, Y => n947);
   U282 : XNOR2X1 port map( A => n171, B => n74, Y => SUMB_10_3_port);
   U283 : XOR2X1 port map( A => CARRYB_9_3_port, B => n577, Y => n171);
   U284 : XNOR2X1 port map( A => n172, B => SUMB_8_10_port, Y => SUMB_9_9_port)
                           ;
   U285 : XNOR2X1 port map( A => ab_9_9_port, B => CARRYB_8_9_port, Y => n172);
   U286 : INVX2 port map( A => n430, Y => n252);
   U287 : NAND2X1 port map( A => ab_1_11_port, B => ab_0_12_port, Y => n174);
   U288 : XOR2X1 port map( A => A(15), B => B(15), Y => n175);
   U289 : XOR2X1 port map( A => n113, B => n175, Y => A1_13_port);
   U290 : NAND2X1 port map( A => SUMB_15_0_port, B => A(15), Y => n176);
   U291 : NAND2X1 port map( A => SUMB_15_0_port, B => B(15), Y => n177);
   U292 : NAND2X1 port map( A => A(15), B => B(15), Y => n178);
   U293 : NAND3X1 port map( A => n178, B => n177, C => n176, Y => A2_14_port);
   U294 : NAND2X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, Y => n928);
   U295 : AND2X1 port map( A => SUMB_15_4_port, B => CARRYB_15_3_port, Y => 
                           n1017);
   U296 : XNOR2X1 port map( A => n235, B => n179, Y => SUMB_8_5_port);
   U297 : XOR2X1 port map( A => CARRYB_7_5_port, B => ab_8_5_port, Y => n179);
   U298 : XOR2X1 port map( A => SUMB_12_8_port, B => n180, Y => SUMB_13_7_port)
                           ;
   U299 : XOR2X1 port map( A => ab_13_7_port, B => CARRYB_12_7_port, Y => n180)
                           ;
   U300 : XOR2X1 port map( A => n181, B => n356, Y => SUMB_3_12_port);
   U301 : XNOR2X1 port map( A => CARRYB_2_12_port, B => ab_3_12_port, Y => n181
                           );
   U302 : INVX2 port map( A => SUMB_13_3_port, Y => n433);
   U303 : XOR2X1 port map( A => n182, B => n68, Y => SUMB_3_9_port);
   U304 : NAND2X1 port map( A => n260, B => n261, Y => n183);
   U305 : NAND3X1 port map( A => n384, B => n383, C => n385, Y => n184);
   U306 : AND2X2 port map( A => ab_0_11_port, B => ab_1_10_port, Y => n185);
   U307 : NAND2X1 port map( A => SUMB_1_13_port, B => n388, Y => n187);
   U308 : NAND2X1 port map( A => SUMB_1_13_port, B => ab_2_12_port, Y => n188);
   U309 : NAND2X1 port map( A => n388, B => ab_2_12_port, Y => n189);
   U310 : NAND3X1 port map( A => n189, B => n187, C => n188, Y => 
                           CARRYB_2_12_port);
   U311 : XNOR2X1 port map( A => n190, B => SUMB_4_12_port, Y => SUMB_5_11_port
                           );
   U312 : XOR2X1 port map( A => n831, B => ab_5_11_port, Y => n190);
   U313 : XOR2X1 port map( A => ab_4_14_port, B => ab_3_15_port, Y => n191);
   U314 : XOR2X1 port map( A => CARRYB_3_14_port, B => n191, Y => 
                           SUMB_4_14_port);
   U315 : NAND2X1 port map( A => CARRYB_3_14_port, B => ab_4_14_port, Y => n192
                           );
   U316 : NAND2X1 port map( A => CARRYB_3_14_port, B => ab_3_15_port, Y => n193
                           );
   U317 : NAND2X1 port map( A => ab_4_14_port, B => ab_3_15_port, Y => n194);
   U318 : NAND3X1 port map( A => n193, B => n192, C => n194, Y => 
                           CARRYB_4_14_port);
   U319 : AND2X2 port map( A => ab_0_15_port, B => ab_1_14_port, Y => n195);
   U320 : AND2X2 port map( A => ab_0_15_port, B => ab_1_14_port, Y => n196);
   U321 : XNOR2X1 port map( A => n197, B => SUMB_10_11_port, Y => n374);
   U322 : XOR2X1 port map( A => SUMB_15_7_port, B => CARRYB_15_6_port, Y => 
                           A1_20_port);
   U323 : NAND2X1 port map( A => ab_4_10_port, B => n834, Y => n198);
   U324 : INVX2 port map( A => n833, Y => n834);
   U325 : XNOR2X1 port map( A => n199, B => SUMB_9_12_port, Y => 
                           SUMB_10_11_port);
   U326 : XNOR2X1 port map( A => CARRYB_9_11_port, B => ab_10_11_port, Y => 
                           n199);
   U327 : XOR2X1 port map( A => n227, B => n431, Y => n200);
   U328 : NAND3X1 port map( A => n786, B => n788, C => n27, Y => n201);
   U329 : INVX2 port map( A => SUMB_11_4_port, Y => n431);
   U330 : XNOR2X1 port map( A => n202, B => SUMB_3_8_port, Y => SUMB_4_7_port);
   U331 : XNOR2X1 port map( A => n947, B => n680, Y => n202);
   U332 : NAND2X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, Y => n203);
   U333 : BUFX2 port map( A => n865, Y => n204);
   U334 : BUFX2 port map( A => SUMB_2_2_port, Y => n205);
   U335 : NAND2X1 port map( A => n447, B => n446, Y => n206);
   U336 : XNOR2X1 port map( A => n207, B => SUMB_2_9_port, Y => SUMB_3_8_port);
   U337 : XNOR2X1 port map( A => CARRYB_2_8_port, B => ab_3_8_port, Y => n207);
   U338 : INVX2 port map( A => SUMB_7_7_port, Y => n217);
   U339 : XNOR2X1 port map( A => n208, B => n138, Y => n212);
   U340 : XOR2X1 port map( A => n225, B => n209, Y => SUMB_10_9_port);
   U341 : INVX2 port map( A => SUMB_9_10_port, Y => n209);
   U342 : AND2X2 port map( A => ab_0_7_port, B => ab_1_6_port, Y => n210);
   U343 : XNOR2X1 port map( A => n212, B => n254, Y => SUMB_4_6_port);
   U344 : XOR2X1 port map( A => CARRYB_14_4_port, B => ab_15_4_port, Y => n309)
                           ;
   U345 : XOR2X1 port map( A => CARRYB_4_10_port, B => n213, Y => n214);
   U346 : XNOR2X1 port map( A => n214, B => n267, Y => SUMB_5_10_port);
   U347 : XOR2X1 port map( A => n215, B => n222, Y => SUMB_3_6_port);
   U348 : XNOR2X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, Y => n215);
   U349 : XOR2X1 port map( A => n216, B => n272, Y => SUMB_2_10_port);
   U350 : INVX1 port map( A => SUMB_1_11_port, Y => n216);
   U351 : NAND3X1 port map( A => n499, B => n500, C => n501, Y => n219);
   U352 : NAND3X1 port map( A => n817, B => n818, C => n819, Y => n220);
   U353 : NAND3X1 port map( A => n644, B => n646, C => n645, Y => n221);
   U354 : INVX1 port map( A => SUMB_2_7_port, Y => n222);
   U355 : XNOR2X1 port map( A => n976, B => n223, Y => SUMB_2_6_port);
   U356 : INVX1 port map( A => SUMB_1_7_port, Y => n223);
   U357 : XNOR2X1 port map( A => ab_10_9_port, B => CARRYB_9_9_port, Y => n225)
                           ;
   U358 : XNOR2X1 port map( A => n226, B => SUMB_8_11_port, Y => SUMB_9_10_port
                           );
   U359 : XNOR2X1 port map( A => CARRYB_8_10_port, B => ab_9_10_port, Y => n226
                           );
   U360 : XOR2X1 port map( A => n227, B => n431, Y => SUMB_12_3_port);
   U361 : NAND3X1 port map( A => n884, B => n885, C => n886, Y => n229);
   U362 : AND2X1 port map( A => SUMB_15_5_port, B => CARRYB_15_4_port, Y => 
                           n1018);
   U363 : XNOR2X1 port map( A => n274, B => n230, Y => SUMB_3_7_port);
   U364 : XOR2X1 port map( A => CARRYB_2_7_port, B => ab_3_7_port, Y => n230);
   U365 : BUFX4 port map( A => SUMB_6_5_port, Y => n575);
   U366 : BUFX2 port map( A => CARRYB_10_5_port, Y => n231);
   U367 : NAND3X1 port map( A => n461, B => n462, C => n460, Y => n232);
   U368 : XOR2X1 port map( A => n233, B => n55, Y => SUMB_4_8_port);
   U369 : XNOR2X1 port map( A => n913, B => ab_4_8_port, Y => n233);
   U370 : XOR2X1 port map( A => CARRYB_6_9_port, B => n234, Y => n421);
   U371 : NAND2X1 port map( A => ab_10_1_port, B => n1026, Y => n236);
   U372 : BUFX2 port map( A => SUMB_3_5_port, Y => n237);
   U373 : XNOR2X1 port map( A => ab_5_12_port, B => n829, Y => n503);
   U374 : INVX2 port map( A => n829, Y => n830);
   U375 : NAND3X1 port map( A => n868, B => n870, C => n869, Y => n238);
   U376 : XNOR2X1 port map( A => n239, B => SUMB_2_6_port, Y => SUMB_3_5_port);
   U377 : XOR2X1 port map( A => ab_3_5_port, B => n985, Y => n239);
   U378 : XOR2X1 port map( A => n240, B => n241, Y => SUMB_11_4_port);
   U379 : XOR2X1 port map( A => n281, B => n519, Y => n241);
   U380 : NAND2X1 port map( A => n790, B => n98, Y => n946);
   U381 : BUFX2 port map( A => n750, Y => n242);
   U382 : INVX1 port map( A => CARRYB_4_2_port, Y => n573);
   U383 : INVX1 port map( A => ab_3_13_port, Y => n244);
   U384 : XNOR2X1 port map( A => n243, B => SUMB_7_11_port, Y => SUMB_8_10_port
                           );
   U385 : XNOR2X1 port map( A => ab_8_10_port, B => CARRYB_7_10_port, Y => n243
                           );
   U386 : XNOR2X1 port map( A => n244, B => CARRYB_2_13_port, Y => n874);
   U387 : INVX2 port map( A => SUMB_8_4_port, Y => n329);
   U388 : BUFX2 port map( A => SUMB_15_3_port, Y => n245);
   U389 : XNOR2X1 port map( A => n246, B => SUMB_14_7_port, Y => SUMB_15_6_port
                           );
   U390 : XOR2X1 port map( A => CARRYB_14_6_port, B => n540, Y => n246);
   U391 : NAND2X1 port map( A => n379, B => n99, Y => n594);
   U392 : INVX2 port map( A => CARRYB_11_1_port, Y => n666);
   U393 : XNOR2X1 port map( A => n247, B => SUMB_10_10_port, Y => 
                           SUMB_11_9_port);
   U394 : XNOR2X1 port map( A => ab_11_9_port, B => CARRYB_10_9_port, Y => n247
                           );
   U395 : XOR2X1 port map( A => n248, B => n527, Y => SUMB_5_4_port);
   U396 : XNOR2X1 port map( A => CARRYB_4_4_port, B => ab_5_4_port, Y => n248);
   U397 : INVX1 port map( A => B(7), Y => n1046);
   U398 : XNOR2X1 port map( A => n249, B => n722, Y => SUMB_2_8_port);
   U399 : XOR2X1 port map( A => ab_2_8_port, B => n440, Y => n249);
   U400 : INVX2 port map( A => CARRYB_6_11_port, Y => n250);
   U401 : INVX4 port map( A => n250, Y => n251);
   U402 : XNOR2X1 port map( A => n253, B => n262, Y => SUMB_2_7_port);
   U403 : XOR2X1 port map( A => ab_2_7_port, B => n270, Y => n253);
   U404 : INVX1 port map( A => n839, Y => n840);
   U405 : INVX2 port map( A => CARRYB_15_0_port, Y => n749);
   U406 : NAND2X1 port map( A => SUMB_14_3_port, B => n201, Y => n256);
   U407 : NAND2X1 port map( A => SUMB_14_3_port, B => ab_15_2_port, Y => n257);
   U408 : NAND2X1 port map( A => n201, B => ab_15_2_port, Y => n258);
   U409 : NAND3X1 port map( A => n258, B => n256, C => n257, Y => 
                           CARRYB_15_2_port);
   U410 : NAND2X1 port map( A => SUMB_13_4_port, B => n277, Y => n260);
   U411 : NAND2X1 port map( A => n63, B => n259, Y => n261);
   U412 : NAND2X1 port map( A => n260, B => n261, Y => SUMB_14_3_port);
   U413 : INVX1 port map( A => SUMB_13_4_port, Y => n259);
   U414 : BUFX2 port map( A => SUMB_1_8_port, Y => n262);
   U415 : NAND3X1 port map( A => n895, B => n897, C => n16, Y => n263);
   U416 : BUFX2 port map( A => SUMB_9_2_port, Y => n264);
   U417 : NAND3X1 port map( A => n795, B => n796, C => n794, Y => n265);
   U418 : NAND3X1 port map( A => n951, B => n952, C => n953, Y => n266);
   U419 : BUFX2 port map( A => SUMB_4_11_port, Y => n267);
   U420 : NAND3X1 port map( A => n811, B => n812, C => n813, Y => n268);
   U421 : NAND3X1 port map( A => n647, B => n648, C => n649, Y => n269);
   U422 : NAND2X1 port map( A => ab_1_7_port, B => ab_0_8_port, Y => n270);
   U423 : INVX1 port map( A => n985, Y => n986);
   U424 : XOR2X1 port map( A => n1024, B => ab_2_10_port, Y => n272);
   U425 : INVX1 port map( A => CARRYB_6_9_port, Y => n839);
   U426 : XNOR2X1 port map( A => n273, B => SUMB_9_8_port, Y => SUMB_10_7_port)
                           ;
   U427 : INVX1 port map( A => SUMB_2_8_port, Y => n274);
   U428 : XNOR2X1 port map( A => n956, B => n275, Y => SUMB_9_6_port);
   U429 : INVX1 port map( A => SUMB_8_7_port, Y => n275);
   U430 : XOR2X1 port map( A => n678, B => n474, Y => n277);
   U431 : BUFX2 port map( A => SUMB_3_6_port, Y => n278);
   U432 : BUFX2 port map( A => SUMB_10_2_port, Y => n279);
   U433 : INVX2 port map( A => SUMB_3_10_port, Y => n314);
   U434 : BUFX2 port map( A => n740, Y => n280);
   U435 : XNOR2X1 port map( A => n281, B => n519, Y => SUMB_10_5_port);
   U436 : XOR2X1 port map( A => CARRYB_6_13_port, B => ab_7_13_port, Y => n282)
                           ;
   U437 : XOR2X1 port map( A => n282, B => SUMB_6_14_port, Y => SUMB_7_13_port)
                           ;
   U438 : NAND2X1 port map( A => SUMB_6_14_port, B => CARRYB_6_13_port, Y => 
                           n283);
   U439 : NAND2X1 port map( A => SUMB_6_14_port, B => ab_7_13_port, Y => n284);
   U440 : NAND2X1 port map( A => CARRYB_6_13_port, B => ab_7_13_port, Y => n285
                           );
   U441 : NAND3X1 port map( A => n284, B => n283, C => n285, Y => 
                           CARRYB_7_13_port);
   U442 : XOR2X1 port map( A => ab_5_15_port, B => ab_6_14_port, Y => n286);
   U443 : XOR2X1 port map( A => CARRYB_5_14_port, B => n286, Y => 
                           SUMB_6_14_port);
   U444 : NAND2X1 port map( A => CARRYB_5_14_port, B => ab_5_15_port, Y => n287
                           );
   U445 : NAND2X1 port map( A => CARRYB_5_14_port, B => ab_6_14_port, Y => n288
                           );
   U446 : NAND2X1 port map( A => ab_5_15_port, B => ab_6_14_port, Y => n289);
   U447 : NAND3X1 port map( A => n288, B => n287, C => n289, Y => 
                           CARRYB_6_14_port);
   U448 : XOR2X1 port map( A => ab_9_13_port, B => CARRYB_8_13_port, Y => n290)
                           ;
   U449 : XOR2X1 port map( A => n290, B => SUMB_8_14_port, Y => SUMB_9_13_port)
                           ;
   U450 : XOR2X1 port map( A => ab_10_12_port, B => CARRYB_9_12_port, Y => n291
                           );
   U451 : XOR2X1 port map( A => n291, B => SUMB_9_13_port, Y => SUMB_10_12_port
                           );
   U452 : NAND2X1 port map( A => ab_9_13_port, B => CARRYB_8_13_port, Y => n292
                           );
   U453 : NAND2X1 port map( A => ab_9_13_port, B => SUMB_8_14_port, Y => n293);
   U454 : NAND2X1 port map( A => CARRYB_8_13_port, B => SUMB_8_14_port, Y => 
                           n294);
   U455 : NAND3X1 port map( A => n292, B => n293, C => n294, Y => 
                           CARRYB_9_13_port);
   U456 : NAND2X1 port map( A => ab_10_12_port, B => CARRYB_9_12_port, Y => 
                           n295);
   U457 : NAND2X1 port map( A => ab_10_12_port, B => SUMB_9_13_port, Y => n296)
                           ;
   U458 : NAND2X1 port map( A => CARRYB_9_12_port, B => SUMB_9_13_port, Y => 
                           n297);
   U459 : NAND3X1 port map( A => n295, B => n296, C => n297, Y => 
                           CARRYB_10_12_port);
   U460 : BUFX2 port map( A => A(0), Y => n298);
   U461 : XOR2X1 port map( A => SUMB_1_5_port, B => ab_2_4_port, Y => n299);
   U462 : XOR2X1 port map( A => n97, B => n299, Y => SUMB_2_4_port);
   U463 : NAND2X1 port map( A => SUMB_1_5_port, B => n97, Y => n300);
   U464 : NAND2X1 port map( A => n97, B => ab_2_4_port, Y => n301);
   U465 : NAND2X1 port map( A => SUMB_1_5_port, B => ab_2_4_port, Y => n302);
   U466 : NAND3X1 port map( A => n301, B => n300, C => n302, Y => 
                           CARRYB_2_4_port);
   U467 : BUFX2 port map( A => SUMB_4_3_port, Y => n303);
   U468 : INVX4 port map( A => A(3), Y => n1066);
   U469 : NAND2X1 port map( A => SUMB_4_10_port, B => CARRYB_4_9_port, Y => 
                           n304);
   U470 : NAND2X1 port map( A => SUMB_4_10_port, B => ab_5_9_port, Y => n305);
   U471 : NAND2X1 port map( A => CARRYB_4_9_port, B => ab_5_9_port, Y => n306);
   U472 : NAND3X1 port map( A => n306, B => n305, C => n304, Y => 
                           CARRYB_5_9_port);
   U473 : NAND3X1 port map( A => n871, B => n51, C => n117, Y => n307);
   U474 : NAND3X1 port map( A => n131, B => n242, C => n752, Y => n308);
   U475 : XOR2X1 port map( A => n309, B => SUMB_14_5_port, Y => SUMB_15_4_port)
                           ;
   U476 : NAND2X1 port map( A => SUMB_14_5_port, B => n129, Y => n310);
   U477 : NAND2X1 port map( A => SUMB_14_5_port, B => ab_15_4_port, Y => n311);
   U478 : NAND2X1 port map( A => n129, B => ab_15_4_port, Y => n312);
   U479 : NAND3X1 port map( A => n311, B => n310, C => n312, Y => 
                           CARRYB_15_4_port);
   U480 : NAND3X1 port map( A => n805, B => n806, C => n807, Y => n313);
   U481 : XNOR2X1 port map( A => n315, B => n126, Y => SUMB_10_2_port);
   U482 : XOR2X1 port map( A => CARRYB_9_2_port, B => n731, Y => n315);
   U483 : NAND3X1 port map( A => n847, B => n848, C => n849, Y => n316);
   U484 : NAND3X1 port map( A => n933, B => n931, C => n932, Y => n317);
   U485 : NAND3X1 port map( A => n915, B => n916, C => n917, Y => n318);
   U486 : XOR2X1 port map( A => n677, B => n319, Y => SUMB_9_2_port);
   U487 : INVX1 port map( A => SUMB_8_3_port, Y => n319);
   U488 : INVX1 port map( A => CARRYB_3_10_port, Y => n833);
   U489 : XNOR2X1 port map( A => n320, B => n136, Y => SUMB_13_4_port);
   U490 : XOR2X1 port map( A => SUMB_12_5_port, B => n590, Y => n320);
   U491 : AND2X2 port map( A => n139, B => n245, Y => n1016);
   U492 : NAND3X1 port map( A => n965, B => n963, C => n964, Y => n321);
   U493 : NAND3X1 port map( A => n856, B => n858, C => n857, Y => n322);
   U494 : NAND3X1 port map( A => n583, B => n584, C => n582, Y => n323);
   U495 : NAND3X1 port map( A => n706, B => n708, C => n707, Y => n324);
   U496 : NAND3X1 port map( A => n198, B => n816, C => n815, Y => n325);
   U497 : NAND3X1 port map( A => n888, B => n890, C => n889, Y => n326);
   U498 : NAND3X1 port map( A => n808, B => n809, C => n810, Y => n327);
   U499 : NAND3X1 port map( A => n465, B => n170, C => n467, Y => n328);
   U500 : XOR2X1 port map( A => n724, B => n329, Y => SUMB_9_3_port);
   U501 : XOR2X1 port map( A => CARRYB_10_8_port, B => ab_11_8_port, Y => n330)
                           ;
   U502 : XOR2X1 port map( A => n330, B => SUMB_10_9_port, Y => SUMB_11_8_port)
                           ;
   U503 : NAND2X1 port map( A => ab_10_9_port, B => n219, Y => n331);
   U504 : NAND2X1 port map( A => SUMB_9_10_port, B => ab_10_9_port, Y => n332);
   U505 : NAND2X1 port map( A => n219, B => SUMB_9_10_port, Y => n333);
   U506 : NAND3X1 port map( A => n331, B => n332, C => n333, Y => 
                           CARRYB_10_9_port);
   U507 : NAND2X1 port map( A => ab_11_8_port, B => n109, Y => n334);
   U508 : NAND2X1 port map( A => SUMB_10_9_port, B => ab_11_8_port, Y => n335);
   U509 : NAND2X1 port map( A => n109, B => SUMB_10_9_port, Y => n336);
   U510 : NAND3X1 port map( A => n334, B => n335, C => n336, Y => 
                           CARRYB_11_8_port);
   U511 : INVX2 port map( A => CARRYB_15_5_port, Y => n510);
   U512 : NAND2X1 port map( A => SUMB_7_7_port, B => n143, Y => n337);
   U513 : NAND2X1 port map( A => SUMB_7_7_port, B => ab_8_6_port, Y => n338);
   U514 : NAND2X1 port map( A => n143, B => ab_8_6_port, Y => n339);
   U515 : NAND3X1 port map( A => n338, B => n337, C => n339, Y => 
                           CARRYB_8_6_port);
   U516 : NAND3X1 port map( A => n4, B => n280, C => n6, Y => n340);
   U517 : NAND3X1 port map( A => n559, B => n558, C => n557, Y => n341);
   U518 : INVX2 port map( A => n831, Y => n832);
   U519 : XOR2X1 port map( A => SUMB_10_1_port, B => ab_11_0_port, Y => n342);
   U520 : XOR2X1 port map( A => CARRYB_10_0_port, B => n342, Y => A1_9_port);
   U521 : NAND2X1 port map( A => CARRYB_10_0_port, B => SUMB_10_1_port, Y => 
                           n343);
   U522 : NAND2X1 port map( A => CARRYB_10_0_port, B => ab_11_0_port, Y => n344
                           );
   U523 : NAND2X1 port map( A => SUMB_10_1_port, B => ab_11_0_port, Y => n345);
   U524 : NAND3X1 port map( A => n344, B => n343, C => n345, Y => 
                           CARRYB_11_0_port);
   U525 : INVX1 port map( A => CARRYB_11_0_port, Y => n866);
   U526 : XNOR2X1 port map( A => n346, B => SUMB_6_11_port, Y => SUMB_7_10_port
                           );
   U527 : XNOR2X1 port map( A => ab_7_10_port, B => CARRYB_6_10_port, Y => n346
                           );
   U528 : INVX2 port map( A => n866, Y => n867);
   U529 : NAND3X1 port map( A => n236, B => n720, C => n721, Y => n347);
   U530 : INVX1 port map( A => n524, Y => n348);
   U531 : NAND3X1 port map( A => n977, B => n978, C => n979, Y => n349);
   U532 : INVX1 port map( A => SUMB_4_4_port, Y => n522);
   U533 : NAND2X1 port map( A => SUMB_4_11_port, B => n325, Y => n350);
   U534 : NAND2X1 port map( A => SUMB_4_11_port, B => ab_5_10_port, Y => n351);
   U535 : NAND2X1 port map( A => n325, B => ab_5_10_port, Y => n352);
   U536 : NAND3X1 port map( A => n351, B => n350, C => n352, Y => 
                           CARRYB_5_10_port);
   U537 : XOR2X1 port map( A => n354, B => n353, Y => SUMB_6_3_port);
   U538 : XNOR2X1 port map( A => n142, B => ab_6_3_port, Y => n353);
   U539 : INVX1 port map( A => SUMB_5_4_port, Y => n354);
   U540 : XNOR2X1 port map( A => n426, B => n264, Y => SUMB_10_1_port);
   U541 : INVX1 port map( A => n1056, Y => n1084);
   U542 : XNOR2X1 port map( A => n357, B => SUMB_9_9_port, Y => SUMB_10_8_port)
                           ;
   U543 : XOR2X1 port map( A => ab_6_13_port, B => CARRYB_5_13_port, Y => n358)
                           ;
   U544 : XOR2X1 port map( A => n358, B => SUMB_5_14_port, Y => SUMB_6_13_port)
                           ;
   U545 : XOR2X1 port map( A => ab_7_12_port, B => CARRYB_6_12_port, Y => n359)
                           ;
   U546 : XOR2X1 port map( A => n359, B => SUMB_6_13_port, Y => SUMB_7_12_port)
                           ;
   U547 : NAND2X1 port map( A => ab_6_13_port, B => CARRYB_5_13_port, Y => n360
                           );
   U548 : NAND2X1 port map( A => ab_6_13_port, B => SUMB_5_14_port, Y => n361);
   U549 : NAND2X1 port map( A => CARRYB_5_13_port, B => SUMB_5_14_port, Y => 
                           n362);
   U550 : NAND3X1 port map( A => n360, B => n361, C => n362, Y => 
                           CARRYB_6_13_port);
   U551 : NAND2X1 port map( A => ab_7_12_port, B => CARRYB_6_12_port, Y => n363
                           );
   U552 : NAND2X1 port map( A => ab_7_12_port, B => SUMB_6_13_port, Y => n364);
   U553 : NAND2X1 port map( A => CARRYB_6_12_port, B => SUMB_6_13_port, Y => 
                           n365);
   U554 : NAND3X1 port map( A => n363, B => n364, C => n365, Y => 
                           CARRYB_7_12_port);
   U555 : XOR2X1 port map( A => CARRYB_12_8_port, B => ab_13_8_port, Y => n366)
                           ;
   U556 : XOR2X1 port map( A => SUMB_12_9_port, B => n366, Y => SUMB_13_8_port)
                           ;
   U557 : NAND2X1 port map( A => SUMB_12_9_port, B => CARRYB_12_8_port, Y => 
                           n367);
   U558 : NAND2X1 port map( A => SUMB_12_9_port, B => ab_13_8_port, Y => n368);
   U559 : NAND2X1 port map( A => CARRYB_12_8_port, B => ab_13_8_port, Y => n369
                           );
   U560 : NAND3X1 port map( A => n368, B => n367, C => n369, Y => 
                           CARRYB_13_8_port);
   U561 : XOR2X1 port map( A => ab_10_10_port, B => CARRYB_9_10_port, Y => n370
                           );
   U562 : XOR2X1 port map( A => n370, B => SUMB_9_11_port, Y => SUMB_10_10_port
                           );
   U563 : NAND2X1 port map( A => ab_10_10_port, B => CARRYB_9_10_port, Y => 
                           n371);
   U564 : NAND2X1 port map( A => ab_10_10_port, B => SUMB_9_11_port, Y => n372)
                           ;
   U565 : NAND2X1 port map( A => CARRYB_9_10_port, B => SUMB_9_11_port, Y => 
                           n373);
   U566 : NAND3X1 port map( A => n371, B => n372, C => n373, Y => 
                           CARRYB_10_10_port);
   U567 : XOR2X1 port map( A => n374, B => CARRYB_10_10_port, Y => 
                           SUMB_11_10_port);
   U568 : NAND2X1 port map( A => ab_11_10_port, B => n19, Y => n375);
   U569 : NAND2X1 port map( A => ab_11_10_port, B => CARRYB_10_10_port, Y => 
                           n376);
   U570 : NAND2X1 port map( A => n19, B => CARRYB_10_10_port, Y => n377);
   U571 : NAND3X1 port map( A => n375, B => n376, C => n377, Y => 
                           CARRYB_11_10_port);
   U572 : XNOR2X1 port map( A => n435, B => SUMB_8_9_port, Y => SUMB_9_8_port);
   U573 : XOR2X1 port map( A => n347, B => ab_11_1_port, Y => n378);
   U574 : XOR2X1 port map( A => n279, B => n378, Y => SUMB_11_1_port);
   U575 : NAND2X1 port map( A => CARRYB_10_1_port, B => SUMB_10_2_port, Y => 
                           n379);
   U576 : NAND2X1 port map( A => SUMB_10_2_port, B => ab_11_1_port, Y => n380);
   U577 : NAND2X1 port map( A => CARRYB_10_1_port, B => ab_11_1_port, Y => n381
                           );
   U578 : NAND3X1 port map( A => n380, B => n379, C => n381, Y => 
                           CARRYB_11_1_port);
   U579 : INVX1 port map( A => n1045, Y => n1088);
   U580 : XNOR2X1 port map( A => n382, B => SUMB_4_6_port, Y => SUMB_5_5_port);
   U581 : XOR2X1 port map( A => CARRYB_4_5_port, B => n434, Y => n382);
   U582 : NAND2X1 port map( A => SUMB_1_12_port, B => n186, Y => n383);
   U583 : NAND2X1 port map( A => SUMB_1_12_port, B => n106, Y => n384);
   U584 : NAND2X1 port map( A => n186, B => n106, Y => n385);
   U585 : INVX4 port map( A => B(12), Y => n1055);
   U586 : XOR2X1 port map( A => n386, B => n387, Y => SUMB_13_3_port);
   U587 : AND2X2 port map( A => ab_0_13_port, B => ab_1_12_port, Y => n388);
   U588 : NAND3X1 port map( A => n709, B => n710, C => n711, Y => n389);
   U589 : NAND3X1 port map( A => n457, B => n456, C => n458, Y => n390);
   U590 : NAND3X1 port map( A => n512, B => n513, C => n514, Y => n391);
   U591 : XNOR2X1 port map( A => ab_0_10_port, B => n392, Y => SUMB_1_9_port);
   U592 : NAND2X1 port map( A => n983, B => n1050, Y => n392);
   U593 : NAND3X1 port map( A => n565, B => n563, C => n564, Y => n393);
   U594 : NAND3X1 port map( A => n898, B => n900, C => n57, Y => n395);
   U595 : NAND3X1 port map( A => n934, B => n935, C => n936, Y => n396);
   U596 : INVX1 port map( A => CARRYB_10_7_port, Y => n657);
   U597 : XOR2X1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, Y => n398)
                           ;
   U598 : XOR2X1 port map( A => n398, B => SUMB_8_13_port, Y => SUMB_9_12_port)
                           ;
   U599 : NAND2X1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, Y => n399
                           );
   U600 : NAND2X1 port map( A => ab_9_12_port, B => SUMB_8_13_port, Y => n400);
   U601 : NAND2X1 port map( A => CARRYB_8_12_port, B => SUMB_8_13_port, Y => 
                           n401);
   U602 : NAND3X1 port map( A => n399, B => n400, C => n401, Y => 
                           CARRYB_9_12_port);
   U603 : NAND2X1 port map( A => ab_10_11_port, B => CARRYB_9_11_port, Y => 
                           n402);
   U604 : NAND2X1 port map( A => ab_10_11_port, B => SUMB_9_12_port, Y => n403)
                           ;
   U605 : NAND2X1 port map( A => CARRYB_9_11_port, B => SUMB_9_12_port, Y => 
                           n404);
   U606 : NAND3X1 port map( A => n402, B => n403, C => n404, Y => 
                           CARRYB_10_11_port);
   U607 : XOR2X1 port map( A => ab_5_13_port, B => CARRYB_4_13_port, Y => n405)
                           ;
   U608 : XOR2X1 port map( A => n405, B => SUMB_4_14_port, Y => SUMB_5_13_port)
                           ;
   U609 : NAND2X1 port map( A => ab_5_13_port, B => CARRYB_4_13_port, Y => n406
                           );
   U610 : NAND2X1 port map( A => ab_5_13_port, B => SUMB_4_14_port, Y => n407);
   U611 : NAND2X1 port map( A => CARRYB_4_13_port, B => SUMB_4_14_port, Y => 
                           n408);
   U612 : NAND3X1 port map( A => n406, B => n407, C => n408, Y => 
                           CARRYB_5_13_port);
   U613 : NAND2X1 port map( A => ab_6_12_port, B => CARRYB_5_12_port, Y => n409
                           );
   U614 : NAND2X1 port map( A => ab_6_12_port, B => SUMB_5_13_port, Y => n410);
   U615 : NAND2X1 port map( A => CARRYB_5_12_port, B => SUMB_5_13_port, Y => 
                           n411);
   U616 : NAND3X1 port map( A => n409, B => n410, C => n411, Y => 
                           CARRYB_6_12_port);
   U617 : XNOR2X1 port map( A => n412, B => SUMB_5_11_port, Y => SUMB_6_10_port
                           );
   U618 : XOR2X1 port map( A => ab_6_10_port, B => n837, Y => n412);
   U619 : XOR2X1 port map( A => SUMB_11_1_port, B => ab_12_0_port, Y => n413);
   U620 : XOR2X1 port map( A => n867, B => n413, Y => A1_10_port);
   U621 : NAND2X1 port map( A => CARRYB_11_0_port, B => SUMB_11_1_port, Y => 
                           n414);
   U622 : NAND2X1 port map( A => CARRYB_11_0_port, B => ab_12_0_port, Y => n415
                           );
   U623 : NAND2X1 port map( A => SUMB_11_1_port, B => ab_12_0_port, Y => n416);
   U624 : NAND3X1 port map( A => n415, B => n416, C => n414, Y => 
                           CARRYB_12_0_port);
   U625 : BUFX2 port map( A => SUMB_5_3_port, Y => n417);
   U626 : NAND3X1 port map( A => n864, B => n863, C => n204, Y => n418);
   U627 : NAND3X1 port map( A => n980, B => n982, C => n981, Y => n419);
   U628 : NAND3X1 port map( A => n472, B => n471, C => n473, Y => n420);
   U629 : XNOR2X1 port map( A => n421, B => SUMB_6_10_port, Y => SUMB_7_9_port)
                           ;
   U630 : NAND3X1 port map( A => n960, B => n961, C => n962, Y => n422);
   U631 : NAND2X1 port map( A => ab_7_2_port, B => n5, Y => n423);
   U632 : BUFX2 port map( A => SUMB_2_5_port, Y => n424);
   U633 : XOR2X1 port map( A => n425, B => n660, Y => SUMB_2_5_port);
   U634 : XNOR2X1 port map( A => n439, B => ab_2_5_port, Y => n425);
   U635 : XNOR2X1 port map( A => n1026, B => ab_10_1_port, Y => n426);
   U636 : NAND3X1 port map( A => n203, B => n638, C => n639, Y => n427);
   U637 : NAND3X1 port map( A => n998, B => n997, C => n999, Y => n428);
   U638 : AND2X2 port map( A => n983, B => n1050, Y => n429);
   U639 : INVX2 port map( A => A(1), Y => n1063);
   U640 : AND2X2 port map( A => n252, B => B(8), Y => ab_1_8_port);
   U641 : XOR2X1 port map( A => n432, B => n433, Y => SUMB_14_2_port);
   U642 : INVX1 port map( A => SUMB_7_5_port, Y => n589);
   U643 : INVX2 port map( A => ab_1_15_port, Y => n511);
   U644 : XNOR2X1 port map( A => CARRYB_8_8_port, B => ab_9_8_port, Y => n435);
   U645 : NAND3X1 port map( A => n630, B => n631, C => n632, Y => n436);
   U646 : AND2X2 port map( A => ab_1_7_port, B => ab_0_8_port, Y => n437);
   U647 : AND2X2 port map( A => B(7), B => n983, Y => ab_1_7_port);
   U648 : INVX1 port map( A => SUMB_1_6_port, Y => n660);
   U649 : INVX2 port map( A => B(8), Y => n1048);
   U650 : INVX2 port map( A => n1063, Y => n984);
   U651 : BUFX2 port map( A => SUMB_3_4_port, Y => n438);
   U652 : AND2X2 port map( A => ab_0_6_port, B => ab_1_5_port, Y => n439);
   U653 : AND2X2 port map( A => n984, B => B(2), Y => n1022);
   U654 : AND2X2 port map( A => ab_1_8_port, B => ab_0_9_port, Y => n440);
   U655 : XNOR2X1 port map( A => n420, B => ab_7_4_port, Y => n441);
   U656 : NAND3X1 port map( A => n923, B => n922, C => n921, Y => n442);
   U657 : XNOR2X1 port map( A => n443, B => n424, Y => SUMB_3_4_port);
   U658 : XOR2X1 port map( A => n701, B => ab_3_4_port, Y => n443);
   U659 : NAND2X1 port map( A => SUMB_6_7_port, B => n626, Y => n446);
   U660 : NAND2X1 port map( A => n444, B => n445, Y => n447);
   U661 : NAND2X1 port map( A => n446, B => n447, Y => SUMB_7_6_port);
   U662 : INVX1 port map( A => n626, Y => n444);
   U663 : INVX1 port map( A => SUMB_6_7_port, Y => n445);
   U664 : XNOR2X1 port map( A => CARRYB_11_2_port, B => n448, Y => n702);
   U665 : XOR2X1 port map( A => n449, B => n450, Y => SUMB_1_7_port);
   U666 : NAND2X1 port map( A => n984, B => B(7), Y => n449);
   U667 : OR2X2 port map( A => n1048, B => n1061, Y => n450);
   U668 : INVX2 port map( A => CARRYB_7_3_port, Y => n524);
   U669 : INVX2 port map( A => n1030, Y => n1031);
   U670 : AND2X2 port map( A => B(15), B => n1061, Y => ab_0_15_port);
   U671 : NAND3X1 port map( A => n712, B => n713, C => n714, Y => n451);
   U672 : XNOR2X1 port map( A => n452, B => SUMB_13_8_port, Y => SUMB_14_7_port
                           );
   U673 : XNOR2X1 port map( A => ab_14_7_port, B => CARRYB_13_7_port, Y => n452
                           );
   U674 : XNOR2X1 port map( A => n1008, B => n453, Y => SUMB_7_2_port);
   U675 : NAND3X1 port map( A => n703, B => n704, C => n705, Y => n454);
   U676 : NAND3X1 port map( A => n907, B => n908, C => n909, Y => n455);
   U677 : NAND2X1 port map( A => SUMB_7_9_port, B => CARRYB_7_8_port, Y => n456
                           );
   U678 : NAND2X1 port map( A => CARRYB_7_8_port, B => ab_8_8_port, Y => n457);
   U679 : NAND2X1 port map( A => SUMB_7_9_port, B => ab_8_8_port, Y => n458);
   U680 : NAND3X1 port map( A => n457, B => n456, C => n458, Y => 
                           CARRYB_8_8_port);
   U681 : XOR2X1 port map( A => SUMB_10_6_port, B => ab_11_5_port, Y => n459);
   U682 : XOR2X1 port map( A => n459, B => n231, Y => SUMB_11_5_port);
   U683 : NAND2X1 port map( A => SUMB_10_6_port, B => CARRYB_10_5_port, Y => 
                           n460);
   U684 : NAND2X1 port map( A => CARRYB_10_5_port, B => ab_11_5_port, Y => n461
                           );
   U685 : NAND2X1 port map( A => SUMB_10_6_port, B => ab_11_5_port, Y => n462);
   U686 : NAND3X1 port map( A => n461, B => n462, C => n460, Y => 
                           CARRYB_11_5_port);
   U687 : XOR2X1 port map( A => CARRYB_7_2_port, B => n463, Y => n673);
   U688 : INVX1 port map( A => n1028, Y => n1029);
   U689 : NAND2X1 port map( A => ab_9_8_port, B => n390, Y => n465);
   U690 : NAND2X1 port map( A => ab_9_8_port, B => SUMB_8_9_port, Y => n466);
   U691 : NAND2X1 port map( A => SUMB_8_9_port, B => n390, Y => n467);
   U692 : NAND3X1 port map( A => n465, B => n466, C => n467, Y => 
                           CARRYB_9_8_port);
   U693 : NAND2X1 port map( A => ab_10_7_port, B => n238, Y => n468);
   U694 : NAND2X1 port map( A => ab_10_7_port, B => SUMB_9_8_port, Y => n469);
   U695 : NAND2X1 port map( A => n238, B => SUMB_9_8_port, Y => n470);
   U696 : NAND3X1 port map( A => n468, B => n469, C => n470, Y => 
                           CARRYB_10_7_port);
   U697 : AND2X2 port map( A => B(9), B => n298, Y => ab_0_9_port);
   U698 : NAND2X1 port map( A => SUMB_5_5_port, B => CARRYB_5_4_port, Y => n471
                           );
   U699 : NAND2X1 port map( A => CARRYB_5_4_port, B => ab_6_4_port, Y => n472);
   U700 : NAND2X1 port map( A => SUMB_5_5_port, B => ab_6_4_port, Y => n473);
   U701 : NAND3X1 port map( A => n472, B => n473, C => n471, Y => 
                           CARRYB_6_4_port);
   U702 : XOR2X1 port map( A => n475, B => n278, Y => SUMB_4_5_port);
   U703 : XOR2X1 port map( A => CARRYB_3_5_port, B => ab_4_5_port, Y => n475);
   U704 : BUFX2 port map( A => SUMB_3_3_port, Y => n476);
   U705 : XNOR2X1 port map( A => n987, B => n477, Y => SUMB_3_3_port);
   U706 : INVX1 port map( A => SUMB_2_4_port, Y => n477);
   U707 : XNOR2X1 port map( A => n676, B => n478, Y => SUMB_7_3_port);
   U708 : XOR2X1 port map( A => CARRYB_6_3_port, B => ab_7_3_port, Y => n478);
   U709 : XOR2X1 port map( A => SUMB_8_1_port, B => ab_9_0_port, Y => n479);
   U710 : XOR2X1 port map( A => n479, B => CARRYB_8_0_port, Y => A1_7_port);
   U711 : NAND2X1 port map( A => CARRYB_8_0_port, B => SUMB_8_1_port, Y => n480
                           );
   U712 : NAND2X1 port map( A => CARRYB_8_0_port, B => ab_9_0_port, Y => n481);
   U713 : NAND2X1 port map( A => SUMB_8_1_port, B => ab_9_0_port, Y => n482);
   U714 : NAND3X1 port map( A => n482, B => n480, C => n481, Y => 
                           CARRYB_9_0_port);
   U715 : XOR2X1 port map( A => ab_2_1_port, B => n96, Y => n483);
   U716 : XOR2X1 port map( A => n483, B => SUMB_1_2_port, Y => SUMB_2_1_port);
   U717 : XOR2X1 port map( A => CARRYB_2_0_port, B => ab_3_0_port, Y => n484);
   U718 : XOR2X1 port map( A => n484, B => SUMB_2_1_port, Y => A1_1_port);
   U719 : NAND2X1 port map( A => ab_2_1_port, B => n96, Y => n485);
   U720 : NAND2X1 port map( A => ab_2_1_port, B => SUMB_1_2_port, Y => n486);
   U721 : NAND2X1 port map( A => n96, B => SUMB_1_2_port, Y => n487);
   U722 : NAND3X1 port map( A => n485, B => n486, C => n487, Y => 
                           CARRYB_2_1_port);
   U723 : NAND2X1 port map( A => CARRYB_2_0_port, B => ab_3_0_port, Y => n488);
   U724 : NAND2X1 port map( A => CARRYB_2_0_port, B => SUMB_2_1_port, Y => n489
                           );
   U725 : NAND2X1 port map( A => ab_3_0_port, B => SUMB_2_1_port, Y => n490);
   U726 : NAND3X1 port map( A => n488, B => n489, C => n490, Y => 
                           CARRYB_3_0_port);
   U727 : INVX1 port map( A => n1037, Y => n1092);
   U728 : INVX2 port map( A => SUMB_9_6_port, Y => n519);
   U729 : NAND2X1 port map( A => SUMB_14_4_port, B => n308, Y => n491);
   U730 : NAND2X1 port map( A => SUMB_14_4_port, B => ab_15_3_port, Y => n492);
   U731 : NAND2X1 port map( A => n308, B => ab_15_3_port, Y => n493);
   U732 : NAND3X1 port map( A => n492, B => n491, C => n493, Y => 
                           CARRYB_15_3_port);
   U733 : NAND3X1 port map( A => n957, B => n39, C => n24, Y => n494);
   U734 : NAND3X1 port map( A => n746, B => n748, C => n747, Y => n495);
   U735 : NAND2X1 port map( A => ab_8_10_port, B => n220, Y => n496);
   U736 : NAND2X1 port map( A => ab_8_10_port, B => SUMB_7_11_port, Y => n497);
   U737 : NAND2X1 port map( A => n220, B => SUMB_7_11_port, Y => n498);
   U738 : NAND3X1 port map( A => n496, B => n497, C => n498, Y => 
                           CARRYB_8_10_port);
   U739 : NAND2X1 port map( A => ab_9_9_port, B => n7, Y => n499);
   U740 : NAND2X1 port map( A => SUMB_8_10_port, B => ab_9_9_port, Y => n500);
   U741 : NAND2X1 port map( A => n7, B => SUMB_8_10_port, Y => n501);
   U742 : NAND3X1 port map( A => n499, B => n500, C => n501, Y => 
                           CARRYB_9_9_port);
   U743 : XOR2X1 port map( A => CARRYB_3_13_port, B => ab_4_13_port, Y => n502)
                           ;
   U744 : XOR2X1 port map( A => n502, B => SUMB_3_14_port, Y => SUMB_4_13_port)
                           ;
   U745 : XOR2X1 port map( A => n503, B => n44, Y => SUMB_5_12_port);
   U746 : NAND2X1 port map( A => ab_4_13_port, B => CARRYB_3_13_port, Y => n504
                           );
   U747 : NAND2X1 port map( A => ab_4_13_port, B => SUMB_3_14_port, Y => n505);
   U748 : NAND2X1 port map( A => CARRYB_3_13_port, B => SUMB_3_14_port, Y => 
                           n506);
   U749 : NAND3X1 port map( A => n504, B => n505, C => n506, Y => 
                           CARRYB_4_13_port);
   U750 : NAND2X1 port map( A => ab_5_12_port, B => n830, Y => n507);
   U751 : NAND2X1 port map( A => ab_5_12_port, B => SUMB_4_13_port, Y => n508);
   U752 : NAND2X1 port map( A => n830, B => SUMB_4_13_port, Y => n509);
   U753 : NAND3X1 port map( A => n507, B => n508, C => n509, Y => 
                           CARRYB_5_12_port);
   U754 : XNOR2X1 port map( A => SUMB_15_6_port, B => n510, Y => A1_19_port);
   U755 : NAND2X1 port map( A => ab_2_7_port, B => n437, Y => n512);
   U756 : NAND2X1 port map( A => n437, B => SUMB_1_8_port, Y => n513);
   U757 : NAND2X1 port map( A => ab_2_7_port, B => SUMB_1_8_port, Y => n514);
   U758 : NAND3X1 port map( A => n512, B => n513, C => n514, Y => 
                           CARRYB_2_7_port);
   U759 : NAND2X1 port map( A => ab_3_6_port, B => n349, Y => n515);
   U760 : NAND2X1 port map( A => ab_3_6_port, B => SUMB_2_7_port, Y => n516);
   U761 : NAND2X1 port map( A => SUMB_2_7_port, B => n349, Y => n517);
   U762 : NAND3X1 port map( A => n515, B => n516, C => n517, Y => 
                           CARRYB_3_6_port);
   U763 : XNOR2X1 port map( A => n441, B => n575, Y => n518);
   U764 : XNOR2X1 port map( A => n954, B => n77, Y => SUMB_15_0_port);
   U765 : OR2X2 port map( A => n520, B => n797, Y => n783);
   U766 : INVX1 port map( A => n797, Y => n798);
   U767 : INVX1 port map( A => n1060, Y => n1082);
   U768 : XOR2X1 port map( A => n522, B => n521, Y => SUMB_5_3_port);
   U769 : XNOR2X1 port map( A => n531, B => ab_5_3_port, Y => n521);
   U770 : NAND2X1 port map( A => n523, B => n524, Y => n525);
   U771 : NAND2X1 port map( A => n973, B => n525, Y => n528);
   U772 : INVX1 port map( A => ab_8_3_port, Y => n523);
   U773 : INVX2 port map( A => n835, Y => n836);
   U774 : XNOR2X1 port map( A => n528, B => n518, Y => SUMB_8_3_port);
   U775 : INVX4 port map( A => n1048, Y => n529);
   U776 : INVX4 port map( A => B(14), Y => n1059);
   U777 : INVX1 port map( A => n837, Y => n838);
   U778 : XNOR2X1 port map( A => n530, B => SUMB_7_10_port, Y => SUMB_8_9_port)
                           ;
   U779 : XNOR2X1 port map( A => CARRYB_7_9_port, B => ab_8_9_port, Y => n530);
   U780 : NAND3X1 port map( A => n665, B => n663, C => n664, Y => n531);
   U781 : INVX2 port map( A => SUMB_5_8_port, Y => n742);
   U782 : XNOR2X1 port map( A => n318, B => n532, Y => n924);
   U783 : NAND2X1 port map( A => SUMB_1_11_port, B => n185, Y => n533);
   U784 : NAND2X1 port map( A => SUMB_1_11_port, B => n104, Y => n534);
   U785 : NAND2X1 port map( A => n104, B => n185, Y => n535);
   U786 : NAND3X1 port map( A => n535, B => n533, C => n534, Y => 
                           CARRYB_2_10_port);
   U787 : INVX4 port map( A => n1049, Y => n579);
   U788 : NAND3X1 port map( A => n853, B => n855, C => n854, Y => n536);
   U789 : NAND3X1 port map( A => n928, B => n930, C => n929, Y => n537);
   U790 : BUFX2 port map( A => SUMB_13_1_port, Y => n538);
   U791 : XNOR2X1 port map( A => n539, B => n82, Y => SUMB_4_11_port);
   U792 : XNOR2X1 port map( A => CARRYB_3_11_port, B => ab_4_11_port, Y => n539
                           );
   U793 : XOR2X1 port map( A => n542, B => n541, Y => SUMB_6_9_port);
   U794 : INVX1 port map( A => SUMB_5_10_port, Y => n542);
   U795 : BUFX2 port map( A => CARRYB_12_0_port, Y => n543);
   U796 : BUFX2 port map( A => SUMB_7_2_port, Y => n544);
   U797 : NAND3X1 port map( A => n923, B => n922, C => n921, Y => n545);
   U798 : NAND3X1 port map( A => n850, B => n851, C => n852, Y => n546);
   U799 : XOR2X1 port map( A => n547, B => n137, Y => SUMB_15_1_port);
   U800 : NAND2X1 port map( A => SUMB_14_2_port, B => n321, Y => n548);
   U801 : NAND2X1 port map( A => SUMB_14_2_port, B => ab_15_1_port, Y => n549);
   U802 : NAND2X1 port map( A => n321, B => ab_15_1_port, Y => n550);
   U803 : NAND3X1 port map( A => n550, B => n548, C => n549, Y => 
                           CARRYB_15_1_port);
   U804 : NAND2X1 port map( A => CARRYB_11_3_port, B => ab_12_3_port, Y => n551
                           );
   U805 : NAND2X1 port map( A => SUMB_11_4_port, B => ab_12_3_port, Y => n552);
   U806 : NAND2X1 port map( A => SUMB_11_4_port, B => CARRYB_11_3_port, Y => 
                           n553);
   U807 : NAND3X1 port map( A => n551, B => n552, C => n553, Y => 
                           CARRYB_12_3_port);
   U808 : NAND2X1 port map( A => ab_13_2_port, B => n324, Y => n554);
   U809 : NAND2X1 port map( A => SUMB_12_3_port, B => ab_13_2_port, Y => n555);
   U810 : NAND2X1 port map( A => SUMB_12_3_port, B => n324, Y => n556);
   U811 : NAND3X1 port map( A => n554, B => n555, C => n556, Y => 
                           CARRYB_13_2_port);
   U812 : NAND2X1 port map( A => n69, B => ab_2_9_port, Y => n557);
   U813 : NAND2X1 port map( A => n69, B => SUMB_1_10_port, Y => n558);
   U814 : NAND2X1 port map( A => SUMB_1_10_port, B => ab_2_9_port, Y => n559);
   U815 : NAND3X1 port map( A => n557, B => n559, C => n558, Y => 
                           CARRYB_2_9_port);
   U816 : NAND2X1 port map( A => ab_3_8_port, B => n396, Y => n560);
   U817 : NAND2X1 port map( A => SUMB_2_9_port, B => ab_3_8_port, Y => n561);
   U818 : NAND2X1 port map( A => SUMB_2_9_port, B => n396, Y => n562);
   U819 : NAND3X1 port map( A => n560, B => n561, C => n562, Y => 
                           CARRYB_3_8_port);
   U820 : NAND2X1 port map( A => n206, B => n536, Y => n563);
   U821 : NAND2X1 port map( A => SUMB_7_6_port, B => ab_8_5_port, Y => n564);
   U822 : NAND2X1 port map( A => n536, B => ab_8_5_port, Y => n565);
   U823 : NAND3X1 port map( A => n565, B => n563, C => n564, Y => 
                           CARRYB_8_5_port);
   U824 : NAND2X1 port map( A => n943, B => n945, Y => n566);
   U825 : NAND2X1 port map( A => n944, B => n567, Y => n969);
   U826 : INVX2 port map( A => n566, Y => n567);
   U827 : XNOR2X1 port map( A => n568, B => n237, Y => SUMB_4_4_port);
   U828 : XNOR2X1 port map( A => ab_4_4_port, B => n266, Y => n568);
   U829 : XNOR2X1 port map( A => n569, B => n60, Y => SUMB_3_10_port);
   U830 : XNOR2X1 port map( A => ab_3_10_port, B => CARRYB_2_10_port, Y => n569
                           );
   U831 : XNOR2X1 port map( A => n570, B => SUMB_13_5_port, Y => SUMB_14_4_port
                           );
   U832 : XNOR2X1 port map( A => ab_14_4_port, B => CARRYB_13_4_port, Y => n570
                           );
   U833 : NAND3X1 port map( A => n602, B => n601, C => n8, Y => n571);
   U834 : NAND2X1 port map( A => n572, B => n573, Y => n574);
   U835 : NAND2X1 port map( A => n635, B => n574, Y => n578);
   U836 : INVX1 port map( A => ab_5_2_port, Y => n572);
   U837 : XNOR2X1 port map( A => n576, B => n544, Y => SUMB_8_1_port);
   U838 : XNOR2X1 port map( A => ab_8_1_port, B => n428, Y => n576);
   U839 : XNOR2X1 port map( A => n578, B => n303, Y => SUMB_5_2_port);
   U840 : INVX1 port map( A => n1049, Y => n1050);
   U841 : INVX2 port map( A => B(9), Y => n1049);
   U842 : NAND3X1 port map( A => n918, B => n920, C => n919, Y => n580);
   U843 : NAND3X1 port map( A => n970, B => n971, C => n972, Y => n581);
   U844 : INVX4 port map( A => n1063, Y => n983);
   U845 : NAND2X1 port map( A => SUMB_5_6_port, B => n580, Y => n582);
   U846 : NAND2X1 port map( A => SUMB_5_6_port, B => ab_6_5_port, Y => n583);
   U847 : NAND2X1 port map( A => n580, B => ab_6_5_port, Y => n584);
   U848 : NAND3X1 port map( A => n583, B => n584, C => n582, Y => 
                           CARRYB_6_5_port);
   U849 : NAND2X1 port map( A => ab_9_6_port, B => n586, Y => n587);
   U850 : NAND2X1 port map( A => CARRYB_8_6_port, B => n585, Y => n588);
   U851 : NAND2X1 port map( A => n587, B => n588, Y => n956);
   U852 : INVX1 port map( A => ab_9_6_port, Y => n585);
   U853 : INVX1 port map( A => CARRYB_8_6_port, Y => n586);
   U854 : NAND2X1 port map( A => SUMB_11_7_port, B => CARRYB_11_6_port, Y => 
                           n591);
   U855 : NAND2X1 port map( A => CARRYB_11_6_port, B => ab_12_6_port, Y => n592
                           );
   U856 : NAND2X1 port map( A => SUMB_11_7_port, B => ab_12_6_port, Y => n593);
   U857 : NAND3X1 port map( A => n592, B => n591, C => n593, Y => 
                           CARRYB_12_6_port);
   U858 : NAND2X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, Y => n595);
   U859 : NAND2X1 port map( A => ab_4_4_port, B => SUMB_3_5_port, Y => n596);
   U860 : NAND2X1 port map( A => CARRYB_3_4_port, B => SUMB_3_5_port, Y => n597
                           );
   U861 : NAND3X1 port map( A => n595, B => n596, C => n597, Y => 
                           CARRYB_4_4_port);
   U862 : NAND2X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, Y => n598);
   U863 : NAND2X1 port map( A => ab_5_3_port, B => SUMB_4_4_port, Y => n599);
   U864 : NAND2X1 port map( A => SUMB_4_4_port, B => CARRYB_4_3_port, Y => n600
                           );
   U865 : NAND2X1 port map( A => n419, B => SUMB_3_6_port, Y => n601);
   U866 : NAND2X1 port map( A => SUMB_3_6_port, B => ab_4_5_port, Y => n602);
   U867 : NAND2X1 port map( A => n419, B => ab_4_5_port, Y => n603);
   U868 : NAND3X1 port map( A => n602, B => n603, C => n601, Y => 
                           CARRYB_4_5_port);
   U869 : XOR2X1 port map( A => SUMB_6_1_port, B => ab_7_0_port, Y => n604);
   U870 : XOR2X1 port map( A => n661, B => n604, Y => A1_5_port);
   U871 : NAND2X1 port map( A => n661, B => SUMB_6_1_port, Y => n605);
   U872 : NAND2X1 port map( A => n661, B => ab_7_0_port, Y => n606);
   U873 : NAND2X1 port map( A => SUMB_6_1_port, B => ab_7_0_port, Y => n607);
   U874 : NAND3X1 port map( A => n606, B => n605, C => n607, Y => 
                           CARRYB_7_0_port);
   U875 : XOR2X1 port map( A => SUMB_3_2_port, B => ab_4_1_port, Y => n608);
   U876 : XOR2X1 port map( A => CARRYB_3_1_port, B => n608, Y => SUMB_4_1_port)
                           ;
   U877 : NAND2X1 port map( A => CARRYB_3_1_port, B => SUMB_3_2_port, Y => n609
                           );
   U878 : NAND2X1 port map( A => CARRYB_3_1_port, B => ab_4_1_port, Y => n610);
   U879 : NAND2X1 port map( A => SUMB_3_2_port, B => ab_4_1_port, Y => n611);
   U880 : NAND3X1 port map( A => n610, B => n609, C => n611, Y => 
                           CARRYB_4_1_port);
   U881 : XOR2X1 port map( A => ab_2_2_port, B => n78, Y => n612);
   U882 : XOR2X1 port map( A => n612, B => SUMB_1_3_port, Y => SUMB_2_2_port);
   U883 : XOR2X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, Y => n613);
   U884 : XOR2X1 port map( A => n613, B => n205, Y => SUMB_3_1_port);
   U885 : NAND2X1 port map( A => ab_2_2_port, B => n78, Y => n614);
   U886 : NAND2X1 port map( A => ab_2_2_port, B => SUMB_1_3_port, Y => n615);
   U887 : NAND2X1 port map( A => n78, B => SUMB_1_3_port, Y => n616);
   U888 : NAND3X1 port map( A => n614, B => n615, C => n616, Y => 
                           CARRYB_2_2_port);
   U889 : NAND2X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, Y => n617);
   U890 : NAND2X1 port map( A => ab_3_1_port, B => SUMB_2_2_port, Y => n618);
   U891 : NAND2X1 port map( A => CARRYB_2_1_port, B => SUMB_2_2_port, Y => n619
                           );
   U892 : NAND3X1 port map( A => n617, B => n618, C => n619, Y => 
                           CARRYB_3_1_port);
   U893 : XOR2X1 port map( A => CARRYB_4_1_port, B => ab_5_1_port, Y => n620);
   U894 : XOR2X1 port map( A => n625, B => n620, Y => SUMB_5_1_port);
   U895 : NAND2X1 port map( A => SUMB_4_2_port, B => CARRYB_4_1_port, Y => n621
                           );
   U896 : NAND2X1 port map( A => SUMB_4_2_port, B => ab_5_1_port, Y => n622);
   U897 : NAND2X1 port map( A => CARRYB_4_1_port, B => ab_5_1_port, Y => n623);
   U898 : NAND3X1 port map( A => n622, B => n621, C => n623, Y => 
                           CARRYB_5_1_port);
   U899 : BUFX2 port map( A => SUMB_2_3_port, Y => n624);
   U900 : BUFX2 port map( A => SUMB_4_2_port, Y => n625);
   U901 : XNOR2X1 port map( A => CARRYB_6_6_port, B => ab_7_6_port, Y => n626);
   U902 : NAND2X1 port map( A => CARRYB_4_4_port, B => ab_5_4_port, Y => n627);
   U903 : NAND2X1 port map( A => SUMB_4_5_port, B => CARRYB_4_4_port, Y => n628
                           );
   U904 : NAND2X1 port map( A => SUMB_4_5_port, B => ab_5_4_port, Y => n629);
   U905 : NAND3X1 port map( A => n627, B => n628, C => n629, Y => 
                           CARRYB_5_4_port);
   U906 : NAND2X1 port map( A => ab_6_3_port, B => n56, Y => n630);
   U907 : NAND2X1 port map( A => SUMB_5_4_port, B => ab_6_3_port, Y => n631);
   U908 : NAND2X1 port map( A => SUMB_5_4_port, B => n56, Y => n632);
   U909 : NAND3X1 port map( A => n630, B => n631, C => n632, Y => 
                           CARRYB_6_3_port);
   U910 : NAND3X1 port map( A => n728, B => n729, C => n730, Y => n633);
   U911 : XOR2X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, Y => n634);
   U912 : XOR2X1 port map( A => n634, B => n17, Y => SUMB_6_1_port);
   U913 : NAND2X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, Y => n635);
   U914 : NAND2X1 port map( A => ab_5_2_port, B => SUMB_4_3_port, Y => n636);
   U915 : NAND2X1 port map( A => SUMB_4_3_port, B => CARRYB_4_2_port, Y => n637
                           );
   U916 : NAND3X1 port map( A => n635, B => n637, C => n636, Y => 
                           CARRYB_5_2_port);
   U917 : NAND2X1 port map( A => ab_6_1_port, B => SUMB_5_2_port, Y => n638);
   U918 : NAND2X1 port map( A => CARRYB_5_1_port, B => SUMB_5_2_port, Y => n639
                           );
   U919 : NAND3X1 port map( A => n203, B => n638, C => n639, Y => 
                           CARRYB_6_1_port);
   U920 : INVX2 port map( A => ab_11_7_port, Y => n654);
   U921 : INVX2 port map( A => ab_4_7_port, Y => n680);
   U922 : NAND2X1 port map( A => SUMB_14_6_port, B => CARRYB_14_5_port, Y => 
                           n640);
   U923 : NAND2X1 port map( A => SUMB_14_6_port, B => ab_15_5_port, Y => n641);
   U924 : NAND2X1 port map( A => CARRYB_14_5_port, B => ab_15_5_port, Y => n642
                           );
   U925 : NAND3X1 port map( A => n641, B => n640, C => n642, Y => 
                           CARRYB_15_5_port);
   U926 : XOR2X1 port map( A => ab_14_6_port, B => CARRYB_13_6_port, Y => n643)
                           ;
   U927 : XOR2X1 port map( A => n643, B => SUMB_13_7_port, Y => SUMB_14_6_port)
                           ;
   U928 : NAND2X1 port map( A => ab_13_7_port, B => CARRYB_12_7_port, Y => n644
                           );
   U929 : NAND2X1 port map( A => ab_13_7_port, B => SUMB_12_8_port, Y => n645);
   U930 : NAND2X1 port map( A => CARRYB_12_7_port, B => SUMB_12_8_port, Y => 
                           n646);
   U931 : NAND3X1 port map( A => n644, B => n646, C => n645, Y => 
                           CARRYB_13_7_port);
   U932 : NAND2X1 port map( A => ab_14_6_port, B => CARRYB_13_6_port, Y => n647
                           );
   U933 : NAND2X1 port map( A => SUMB_13_7_port, B => ab_14_6_port, Y => n648);
   U934 : NAND2X1 port map( A => SUMB_13_7_port, B => CARRYB_13_6_port, Y => 
                           n649);
   U935 : NAND3X1 port map( A => n647, B => n648, C => n649, Y => 
                           CARRYB_14_6_port);
   U936 : XOR2X1 port map( A => CARRYB_11_7_port, B => ab_12_7_port, Y => n650)
                           ;
   U937 : XOR2X1 port map( A => SUMB_11_8_port, B => n650, Y => SUMB_12_7_port)
                           ;
   U938 : NAND2X1 port map( A => SUMB_11_8_port, B => n229, Y => n651);
   U939 : NAND2X1 port map( A => SUMB_11_8_port, B => ab_12_7_port, Y => n652);
   U940 : NAND2X1 port map( A => n229, B => ab_12_7_port, Y => n653);
   U941 : NAND3X1 port map( A => n652, B => n651, C => n653, Y => 
                           CARRYB_12_7_port);
   U942 : INVX1 port map( A => n1043, Y => n1089);
   U943 : INVX1 port map( A => n657, Y => n658);
   U944 : INVX4 port map( A => B(5), Y => n1042);
   U945 : BUFX2 port map( A => CARRYB_3_7_port, Y => n655);
   U946 : NAND3X1 port map( A => n940, B => n941, C => n942, Y => n656);
   U947 : INVX2 port map( A => SUMB_7_3_port, Y => n674);
   U948 : NAND3X1 port map( A => n423, B => n1009, C => n1010, Y => n659);
   U949 : INVX4 port map( A => B(6), Y => n1044);
   U950 : OR2X2 port map( A => n464, B => n1028, Y => n703);
   U951 : BUFX4 port map( A => CARRYB_6_0_port, Y => n661);
   U952 : INVX4 port map( A => B(3), Y => n1038);
   U953 : XOR2X1 port map( A => ab_0_5_port, B => ab_1_4_port, Y => 
                           SUMB_1_4_port);
   U954 : XOR2X1 port map( A => CARRYB_3_3_port, B => ab_4_3_port, Y => n662);
   U955 : XOR2X1 port map( A => n438, B => n662, Y => SUMB_4_3_port);
   U956 : NAND2X1 port map( A => SUMB_3_4_port, B => n145, Y => n663);
   U957 : NAND2X1 port map( A => SUMB_3_4_port, B => ab_4_3_port, Y => n664);
   U958 : NAND2X1 port map( A => n145, B => ab_4_3_port, Y => n665);
   U959 : NAND3X1 port map( A => n664, B => n663, C => n665, Y => 
                           CARRYB_4_3_port);
   U960 : XOR2X1 port map( A => n144, B => ab_6_2_port, Y => n667);
   U961 : XOR2X1 port map( A => n417, B => n667, Y => SUMB_6_2_port);
   U962 : NAND2X1 port map( A => CARRYB_5_2_port, B => SUMB_5_3_port, Y => n668
                           );
   U963 : NAND2X1 port map( A => SUMB_5_3_port, B => ab_6_2_port, Y => n669);
   U964 : NAND2X1 port map( A => CARRYB_5_2_port, B => ab_6_2_port, Y => n670);
   U965 : NAND3X1 port map( A => n670, B => n669, C => n668, Y => 
                           CARRYB_6_2_port);
   U966 : NAND2X1 port map( A => n675, B => CARRYB_6_2_port, Y => n671);
   U967 : NAND2X1 port map( A => ab_7_2_port, B => n1027, Y => n672);
   U968 : NAND2X1 port map( A => n671, B => n672, Y => n1008);
   U969 : INVX1 port map( A => ab_7_2_port, Y => n675);
   U970 : XOR2X1 port map( A => n673, B => n674, Y => SUMB_8_2_port);
   U971 : INVX4 port map( A => B(0), Y => n1032);
   U972 : INVX1 port map( A => SUMB_6_4_port, Y => n676);
   U973 : XNOR2X1 port map( A => n633, B => ab_9_2_port, Y => n677);
   U974 : NAND3X1 port map( A => n783, B => n784, C => n785, Y => n678);
   U975 : NAND3X1 port map( A => n842, B => n841, C => n843, Y => n679);
   U976 : XOR2X1 port map( A => ab_4_12_port, B => CARRYB_3_12_port, Y => n681)
                           ;
   U977 : XOR2X1 port map( A => n681, B => n162, Y => SUMB_4_12_port);
   U978 : NAND2X1 port map( A => ab_4_12_port, B => n128, Y => n682);
   U979 : NAND2X1 port map( A => ab_4_12_port, B => SUMB_3_13_port, Y => n683);
   U980 : NAND2X1 port map( A => n128, B => SUMB_3_13_port, Y => n684);
   U981 : NAND3X1 port map( A => n682, B => n683, C => n684, Y => 
                           CARRYB_4_12_port);
   U982 : NAND2X1 port map( A => ab_5_11_port, B => n832, Y => n685);
   U983 : NAND2X1 port map( A => ab_5_11_port, B => SUMB_4_12_port, Y => n686);
   U984 : NAND2X1 port map( A => n832, B => SUMB_4_12_port, Y => n687);
   U985 : NAND3X1 port map( A => n685, B => n686, C => n687, Y => 
                           CARRYB_5_11_port);
   U986 : NAND2X1 port map( A => ab_14_7_port, B => n221, Y => n688);
   U987 : NAND2X1 port map( A => ab_14_7_port, B => SUMB_13_8_port, Y => n689);
   U988 : NAND2X1 port map( A => n221, B => SUMB_13_8_port, Y => n690);
   U989 : NAND3X1 port map( A => n688, B => n689, C => n690, Y => 
                           CARRYB_14_7_port);
   U990 : NAND2X1 port map( A => ab_15_6_port, B => n269, Y => n691);
   U991 : NAND2X1 port map( A => ab_15_6_port, B => SUMB_14_7_port, Y => n692);
   U992 : NAND2X1 port map( A => n269, B => SUMB_14_7_port, Y => n693);
   U993 : NAND3X1 port map( A => n691, B => n692, C => n693, Y => 
                           CARRYB_15_6_port);
   U994 : NAND2X1 port map( A => ab_11_9_port, B => n135, Y => n694);
   U995 : NAND2X1 port map( A => ab_11_9_port, B => SUMB_10_10_port, Y => n695)
                           ;
   U996 : NAND2X1 port map( A => n135, B => SUMB_10_10_port, Y => n696);
   U997 : NAND3X1 port map( A => n694, B => n695, C => n696, Y => 
                           CARRYB_11_9_port);
   U998 : XOR2X1 port map( A => ab_12_9_port, B => SUMB_11_10_port, Y => n697);
   U999 : XOR2X1 port map( A => n697, B => CARRYB_11_9_port, Y => 
                           SUMB_12_9_port);
   U1000 : NAND2X1 port map( A => ab_12_9_port, B => SUMB_11_10_port, Y => n698
                           );
   U1001 : NAND2X1 port map( A => ab_12_9_port, B => CARRYB_11_9_port, Y => 
                           n699);
   U1002 : NAND2X1 port map( A => SUMB_11_10_port, B => CARRYB_11_9_port, Y => 
                           n700);
   U1003 : NAND3X1 port map( A => n698, B => n699, C => n700, Y => 
                           CARRYB_12_9_port);
   U1004 : INVX2 port map( A => CARRYB_2_4_port, Y => n701);
   U1005 : XOR2X1 port map( A => n702, B => SUMB_11_3_port, Y => SUMB_12_2_port
                           );
   U1006 : NAND2X1 port map( A => SUMB_10_4_port, B => ab_11_3_port, Y => n704)
                           ;
   U1007 : NAND2X1 port map( A => n1029, B => SUMB_10_4_port, Y => n705);
   U1008 : NAND3X1 port map( A => n703, B => n705, C => n704, Y => 
                           CARRYB_11_3_port);
   U1009 : NAND2X1 port map( A => n316, B => ab_12_2_port, Y => n706);
   U1010 : NAND2X1 port map( A => SUMB_11_3_port, B => ab_12_2_port, Y => n707)
                           ;
   U1011 : NAND2X1 port map( A => n316, B => SUMB_11_3_port, Y => n708);
   U1012 : NAND3X1 port map( A => n706, B => n707, C => n708, Y => 
                           CARRYB_12_2_port);
   U1013 : NAND2X1 port map( A => ab_3_9_port, B => n341, Y => n709);
   U1014 : NAND2X1 port map( A => SUMB_2_10_port, B => ab_3_9_port, Y => n710);
   U1015 : NAND2X1 port map( A => SUMB_2_10_port, B => n341, Y => n711);
   U1016 : NAND3X1 port map( A => n709, B => n710, C => n711, Y => 
                           CARRYB_3_9_port);
   U1017 : NAND2X1 port map( A => n914, B => ab_4_8_port, Y => n712);
   U1018 : NAND2X1 port map( A => SUMB_3_9_port, B => ab_4_8_port, Y => n713);
   U1019 : NAND2X1 port map( A => SUMB_3_9_port, B => n914, Y => n714);
   U1020 : NAND3X1 port map( A => n712, B => n713, C => n714, Y => 
                           CARRYB_4_8_port);
   U1021 : XOR2X1 port map( A => n715, B => n742, Y => SUMB_6_7_port);
   U1022 : INVX1 port map( A => n1052, Y => n1085);
   U1023 : INVX2 port map( A => SUMB_1_9_port, Y => n722);
   U1024 : NAND2X1 port map( A => ab_9_2_port, B => CARRYB_8_2_port, Y => n716)
                           ;
   U1025 : NAND2X1 port map( A => SUMB_8_3_port, B => ab_9_2_port, Y => n717);
   U1026 : NAND2X1 port map( A => CARRYB_8_2_port, B => SUMB_8_3_port, Y => 
                           n718);
   U1027 : NAND3X1 port map( A => n716, B => n717, C => n718, Y => 
                           CARRYB_9_2_port);
   U1028 : NAND2X1 port map( A => ab_10_1_port, B => n1026, Y => n719);
   U1029 : NAND2X1 port map( A => ab_10_1_port, B => SUMB_9_2_port, Y => n720);
   U1030 : NAND2X1 port map( A => n1026, B => SUMB_9_2_port, Y => n721);
   U1031 : NAND3X1 port map( A => n719, B => n720, C => n721, Y => 
                           CARRYB_10_1_port);
   U1032 : NAND3X1 port map( A => n975, B => n974, C => n18, Y => n723);
   U1033 : NAND2X1 port map( A => n436, B => ab_7_3_port, Y => n725);
   U1034 : NAND2X1 port map( A => SUMB_6_4_port, B => n436, Y => n726);
   U1035 : NAND2X1 port map( A => SUMB_6_4_port, B => ab_7_3_port, Y => n727);
   U1036 : NAND3X1 port map( A => n725, B => n727, C => n726, Y => 
                           CARRYB_7_3_port);
   U1037 : NAND2X1 port map( A => ab_8_2_port, B => n659, Y => n728);
   U1038 : NAND2X1 port map( A => SUMB_7_3_port, B => ab_8_2_port, Y => n729);
   U1039 : NAND2X1 port map( A => n659, B => SUMB_7_3_port, Y => n730);
   U1040 : NAND3X1 port map( A => n728, B => n729, C => n730, Y => 
                           CARRYB_8_2_port);
   U1041 : INVX1 port map( A => n1047, Y => n1087);
   U1042 : XOR2X1 port map( A => SUMB_1_4_port, B => ab_2_3_port, Y => n732);
   U1043 : XOR2X1 port map( A => n732, B => n1021, Y => SUMB_2_3_port);
   U1044 : NAND2X1 port map( A => SUMB_1_4_port, B => n1021, Y => n733);
   U1045 : NAND2X1 port map( A => n1021, B => ab_2_3_port, Y => n734);
   U1046 : NAND2X1 port map( A => SUMB_1_4_port, B => ab_2_3_port, Y => n735);
   U1047 : NAND3X1 port map( A => n734, B => n733, C => n735, Y => 
                           CARRYB_2_3_port);
   U1048 : INVX4 port map( A => A(2), Y => n1064);
   U1049 : NOR2X1 port map( A => n1061, B => n1044, Y => ab_0_6_port);
   U1050 : NAND2X1 port map( A => n263, B => ab_10_5_port, Y => n736);
   U1051 : NAND2X1 port map( A => SUMB_9_6_port, B => ab_10_5_port, Y => n737);
   U1052 : NAND2X1 port map( A => SUMB_9_6_port, B => n263, Y => n738);
   U1053 : NAND3X1 port map( A => n736, B => n737, C => n738, Y => 
                           CARRYB_10_5_port);
   U1054 : NAND2X1 port map( A => n395, B => ab_11_4_port, Y => n739);
   U1055 : NAND2X1 port map( A => SUMB_10_5_port, B => ab_11_4_port, Y => n740)
                           ;
   U1056 : NAND2X1 port map( A => n395, B => SUMB_10_5_port, Y => n741);
   U1057 : NAND3X1 port map( A => n739, B => n740, C => n741, Y => 
                           CARRYB_11_4_port);
   U1058 : NAND2X1 port map( A => n340, B => ab_12_4_port, Y => n743);
   U1059 : NAND2X1 port map( A => ab_12_4_port, B => SUMB_11_5_port, Y => n744)
                           ;
   U1060 : NAND2X1 port map( A => n340, B => SUMB_11_5_port, Y => n745);
   U1061 : NAND3X1 port map( A => n743, B => n744, C => n745, Y => 
                           CARRYB_12_4_port);
   U1062 : NAND2X1 port map( A => SUMB_12_5_port, B => ab_13_4_port, Y => n746)
                           ;
   U1063 : NAND2X1 port map( A => ab_13_4_port, B => CARRYB_12_4_port, Y => 
                           n747);
   U1064 : NAND2X1 port map( A => SUMB_12_5_port, B => CARRYB_12_4_port, Y => 
                           n748);
   U1065 : NAND3X1 port map( A => n746, B => n747, C => n748, Y => 
                           CARRYB_13_4_port);
   U1066 : INVX1 port map( A => n579, Y => n1086);
   U1067 : XNOR2X1 port map( A => SUMB_15_1_port, B => n749, Y => A1_14_port);
   U1068 : NOR2X1 port map( A => n1061, B => n1048, Y => ab_0_8_port);
   U1069 : NAND2X1 port map( A => SUMB_13_4_port, B => CARRYB_13_3_port, Y => 
                           n750);
   U1070 : NAND2X1 port map( A => SUMB_13_4_port, B => ab_14_3_port, Y => n751)
                           ;
   U1071 : NAND2X1 port map( A => n678, B => ab_14_3_port, Y => n752);
   U1072 : NAND3X1 port map( A => n752, B => n751, C => n750, Y => 
                           CARRYB_14_3_port);
   U1073 : NAND2X1 port map( A => ab_3_10_port, B => n134, Y => n753);
   U1074 : NAND2X1 port map( A => SUMB_2_11_port, B => ab_3_10_port, Y => n754)
                           ;
   U1075 : NAND2X1 port map( A => SUMB_2_11_port, B => n134, Y => n755);
   U1076 : NAND3X1 port map( A => n753, B => n754, C => n755, Y => 
                           CARRYB_3_10_port);
   U1077 : NAND2X1 port map( A => ab_4_9_port, B => n389, Y => n756);
   U1078 : NAND2X1 port map( A => SUMB_3_10_port, B => ab_4_9_port, Y => n757);
   U1079 : NAND2X1 port map( A => SUMB_3_10_port, B => n389, Y => n758);
   U1080 : NAND3X1 port map( A => n756, B => n757, C => n758, Y => 
                           CARRYB_4_9_port);
   U1081 : NAND2X1 port map( A => ab_11_6_port, B => n307, Y => n759);
   U1082 : NAND2X1 port map( A => SUMB_10_7_port, B => ab_11_6_port, Y => n760)
                           ;
   U1083 : NAND2X1 port map( A => SUMB_10_7_port, B => n307, Y => n761);
   U1084 : NAND3X1 port map( A => n759, B => n760, C => n761, Y => 
                           CARRYB_11_6_port);
   U1085 : NAND2X1 port map( A => ab_12_5_port, B => n232, Y => n762);
   U1086 : NAND2X1 port map( A => SUMB_11_6_port, B => ab_12_5_port, Y => n763)
                           ;
   U1087 : NAND2X1 port map( A => SUMB_11_6_port, B => n232, Y => n764);
   U1088 : NAND3X1 port map( A => n762, B => n763, C => n764, Y => 
                           CARRYB_12_5_port);
   U1089 : XOR2X1 port map( A => CARRYB_7_11_port, B => ab_8_11_port, Y => n765
                           );
   U1090 : XOR2X1 port map( A => n765, B => SUMB_7_12_port, Y => SUMB_8_11_port
                           );
   U1091 : NAND2X1 port map( A => ab_8_11_port, B => CARRYB_7_11_port, Y => 
                           n766);
   U1092 : NAND2X1 port map( A => ab_8_11_port, B => SUMB_7_12_port, Y => n767)
                           ;
   U1093 : NAND2X1 port map( A => CARRYB_7_11_port, B => SUMB_7_12_port, Y => 
                           n768);
   U1094 : NAND3X1 port map( A => n766, B => n767, C => n768, Y => 
                           CARRYB_8_11_port);
   U1095 : NAND2X1 port map( A => ab_9_10_port, B => n111, Y => n769);
   U1096 : NAND2X1 port map( A => ab_9_10_port, B => SUMB_8_11_port, Y => n770)
                           ;
   U1097 : NAND2X1 port map( A => n111, B => SUMB_8_11_port, Y => n771);
   U1098 : NAND3X1 port map( A => n769, B => n770, C => n771, Y => 
                           CARRYB_9_10_port);
   U1099 : XOR2X1 port map( A => ab_13_6_port, B => CARRYB_12_6_port, Y => n772
                           );
   U1100 : XOR2X1 port map( A => n772, B => SUMB_12_7_port, Y => SUMB_13_6_port
                           );
   U1101 : NAND2X1 port map( A => ab_13_6_port, B => CARRYB_12_6_port, Y => 
                           n773);
   U1102 : NAND2X1 port map( A => SUMB_12_7_port, B => ab_13_6_port, Y => n774)
                           ;
   U1103 : NAND2X1 port map( A => CARRYB_12_6_port, B => SUMB_12_7_port, Y => 
                           n775);
   U1104 : NAND3X1 port map( A => n773, B => n774, C => n775, Y => 
                           CARRYB_13_6_port);
   U1105 : NAND2X1 port map( A => ab_14_5_port, B => n326, Y => n776);
   U1106 : NAND2X1 port map( A => SUMB_13_6_port, B => ab_14_5_port, Y => n777)
                           ;
   U1107 : NAND2X1 port map( A => n326, B => SUMB_13_6_port, Y => n778);
   U1108 : NAND3X1 port map( A => n776, B => n777, C => n778, Y => 
                           CARRYB_14_5_port);
   U1109 : XOR2X1 port map( A => n779, B => SUMB_1_14_port, Y => SUMB_2_13_port
                           );
   U1110 : NAND2X1 port map( A => SUMB_1_14_port, B => CARRYB_1_13_port, Y => 
                           n780);
   U1111 : NAND2X1 port map( A => SUMB_1_14_port, B => ab_2_13_port, Y => n781)
                           ;
   U1112 : NAND2X1 port map( A => CARRYB_1_13_port, B => ab_2_13_port, Y => 
                           n782);
   U1113 : NAND3X1 port map( A => n782, B => n780, C => n781, Y => 
                           CARRYB_2_13_port);
   U1114 : NAND2X1 port map( A => SUMB_12_4_port, B => ab_13_3_port, Y => n784)
                           ;
   U1115 : NAND2X1 port map( A => SUMB_12_4_port, B => n798, Y => n785);
   U1116 : NAND3X1 port map( A => n783, B => n784, C => n785, Y => 
                           CARRYB_13_3_port);
   U1117 : NAND2X1 port map( A => CARRYB_13_2_port, B => ab_14_2_port, Y => 
                           n786);
   U1118 : NAND2X1 port map( A => SUMB_13_3_port, B => ab_14_2_port, Y => n787)
                           ;
   U1119 : NAND2X1 port map( A => SUMB_13_3_port, B => CARRYB_13_2_port, Y => 
                           n788);
   U1120 : NAND3X1 port map( A => n786, B => n787, C => n788, Y => 
                           CARRYB_14_2_port);
   U1121 : NAND2X1 port map( A => SUMB_4_9_port, B => n451, Y => n789);
   U1122 : NAND2X1 port map( A => SUMB_4_9_port, B => ab_5_8_port, Y => n790);
   U1123 : NAND2X1 port map( A => n451, B => ab_5_8_port, Y => n791);
   U1124 : NAND3X1 port map( A => n791, B => n789, C => n790, Y => 
                           CARRYB_5_8_port);
   U1125 : NAND3X1 port map( A => n901, B => n903, C => n902, Y => n792);
   U1126 : XOR2X1 port map( A => n32, B => ab_13_0_port, Y => n793);
   U1127 : XOR2X1 port map( A => n543, B => n793, Y => A1_11_port);
   U1128 : NAND2X1 port map( A => SUMB_12_1_port, B => CARRYB_12_0_port, Y => 
                           n794);
   U1129 : NAND2X1 port map( A => CARRYB_12_0_port, B => ab_13_0_port, Y => 
                           n795);
   U1130 : NAND2X1 port map( A => SUMB_12_1_port, B => ab_13_0_port, Y => n796)
                           ;
   U1131 : NAND3X1 port map( A => n795, B => n796, C => n794, Y => 
                           CARRYB_13_0_port);
   U1132 : INVX2 port map( A => CARRYB_12_3_port, Y => n797);
   U1133 : NAND2X1 port map( A => ab_6_9_port, B => n836, Y => n799);
   U1134 : NAND2X1 port map( A => SUMB_5_10_port, B => ab_6_9_port, Y => n800);
   U1135 : NAND2X1 port map( A => SUMB_5_10_port, B => n836, Y => n801);
   U1136 : NAND3X1 port map( A => n800, B => n799, C => n801, Y => 
                           CARRYB_6_9_port);
   U1137 : NAND2X1 port map( A => ab_7_8_port, B => n656, Y => n802);
   U1138 : NAND2X1 port map( A => ab_7_8_port, B => SUMB_6_9_port, Y => n803);
   U1139 : NAND2X1 port map( A => n656, B => SUMB_6_9_port, Y => n804);
   U1140 : NAND3X1 port map( A => n802, B => n803, C => n804, Y => 
                           CARRYB_7_8_port);
   U1141 : NAND2X1 port map( A => ab_6_10_port, B => n838, Y => n805);
   U1142 : NAND2X1 port map( A => ab_6_10_port, B => SUMB_5_11_port, Y => n806)
                           ;
   U1143 : NAND2X1 port map( A => n838, B => SUMB_5_11_port, Y => n807);
   U1144 : NAND3X1 port map( A => n805, B => n806, C => n807, Y => 
                           CARRYB_6_10_port);
   U1145 : NAND2X1 port map( A => ab_7_9_port, B => n840, Y => n808);
   U1146 : NAND2X1 port map( A => ab_7_9_port, B => SUMB_6_10_port, Y => n809);
   U1147 : NAND2X1 port map( A => n840, B => SUMB_6_10_port, Y => n810);
   U1148 : NAND3X1 port map( A => n808, B => n809, C => n810, Y => 
                           CARRYB_7_9_port);
   U1149 : NAND2X1 port map( A => ab_3_11_port, B => n184, Y => n811);
   U1150 : NAND2X1 port map( A => SUMB_2_12_port, B => ab_3_11_port, Y => n812)
                           ;
   U1151 : NAND2X1 port map( A => SUMB_2_12_port, B => n184, Y => n813);
   U1152 : NAND3X1 port map( A => n811, B => n812, C => n813, Y => 
                           CARRYB_3_11_port);
   U1153 : NAND2X1 port map( A => ab_4_10_port, B => n834, Y => n814);
   U1154 : NAND2X1 port map( A => SUMB_3_11_port, B => ab_4_10_port, Y => n815)
                           ;
   U1155 : NAND2X1 port map( A => SUMB_3_11_port, B => n834, Y => n816);
   U1156 : NAND3X1 port map( A => n814, B => n815, C => n816, Y => 
                           CARRYB_4_10_port);
   U1157 : NAND2X1 port map( A => ab_7_10_port, B => n313, Y => n817);
   U1158 : NAND2X1 port map( A => ab_7_10_port, B => SUMB_6_11_port, Y => n818)
                           ;
   U1159 : NAND2X1 port map( A => n313, B => SUMB_6_11_port, Y => n819);
   U1160 : NAND3X1 port map( A => n817, B => n818, C => n819, Y => 
                           CARRYB_7_10_port);
   U1161 : NAND2X1 port map( A => ab_8_9_port, B => n327, Y => n820);
   U1162 : NAND2X1 port map( A => ab_8_9_port, B => SUMB_7_10_port, Y => n821);
   U1163 : NAND2X1 port map( A => n327, B => SUMB_7_10_port, Y => n822);
   U1164 : NAND3X1 port map( A => n820, B => n821, C => n822, Y => 
                           CARRYB_8_9_port);
   U1165 : NAND2X1 port map( A => ab_3_12_port, B => n116, Y => n823);
   U1166 : NAND2X1 port map( A => SUMB_2_13_port, B => ab_3_12_port, Y => n824)
                           ;
   U1167 : NAND2X1 port map( A => SUMB_2_13_port, B => n116, Y => n825);
   U1168 : NAND3X1 port map( A => n823, B => n824, C => n825, Y => 
                           CARRYB_3_12_port);
   U1169 : NAND2X1 port map( A => ab_4_11_port, B => n268, Y => n826);
   U1170 : NAND2X1 port map( A => SUMB_3_12_port, B => ab_4_11_port, Y => n827)
                           ;
   U1171 : NAND2X1 port map( A => SUMB_3_12_port, B => n268, Y => n828);
   U1172 : NAND3X1 port map( A => n826, B => n827, C => n828, Y => 
                           CARRYB_4_11_port);
   U1173 : INVX2 port map( A => CARRYB_4_12_port, Y => n829);
   U1174 : INVX2 port map( A => CARRYB_4_11_port, Y => n831);
   U1175 : INVX2 port map( A => CARRYB_5_9_port, Y => n835);
   U1176 : INVX2 port map( A => CARRYB_5_10_port, Y => n837);
   U1177 : NAND2X1 port map( A => n165, B => ab_5_7_port, Y => n841);
   U1178 : NAND2X1 port map( A => SUMB_4_8_port, B => ab_5_7_port, Y => n842);
   U1179 : NAND2X1 port map( A => SUMB_4_8_port, B => n165, Y => n843);
   U1180 : NAND3X1 port map( A => n842, B => n841, C => n843, Y => 
                           CARRYB_5_7_port);
   U1181 : NAND2X1 port map( A => ab_6_6_port, B => n537, Y => n844);
   U1182 : NAND2X1 port map( A => SUMB_5_7_port, B => ab_6_6_port, Y => n845);
   U1183 : NAND2X1 port map( A => n537, B => SUMB_5_7_port, Y => n846);
   U1184 : NAND3X1 port map( A => n844, B => n845, C => n846, Y => 
                           CARRYB_6_6_port);
   U1185 : NAND2X1 port map( A => n442, B => ab_11_2_port, Y => n847);
   U1186 : NAND2X1 port map( A => ab_11_2_port, B => SUMB_10_3_port, Y => n848)
                           ;
   U1187 : NAND2X1 port map( A => n442, B => SUMB_10_3_port, Y => n849);
   U1188 : NAND3X1 port map( A => n847, B => n848, C => n849, Y => 
                           CARRYB_11_2_port);
   U1189 : NAND2X1 port map( A => n594, B => ab_12_1_port, Y => n850);
   U1190 : NAND2X1 port map( A => SUMB_11_2_port, B => ab_12_1_port, Y => n851)
                           ;
   U1191 : NAND2X1 port map( A => SUMB_11_2_port, B => n594, Y => n852);
   U1192 : NAND3X1 port map( A => n851, B => n850, C => n852, Y => 
                           CARRYB_12_1_port);
   U1193 : NAND2X1 port map( A => ab_7_5_port, B => n323, Y => n853);
   U1194 : NAND2X1 port map( A => SUMB_6_6_port, B => ab_7_5_port, Y => n854);
   U1195 : NAND2X1 port map( A => SUMB_6_6_port, B => n323, Y => n855);
   U1196 : NAND3X1 port map( A => n853, B => n854, C => n855, Y => 
                           CARRYB_7_5_port);
   U1197 : NAND2X1 port map( A => ab_8_4_port, B => n581, Y => n856);
   U1198 : NAND2X1 port map( A => SUMB_7_5_port, B => ab_8_4_port, Y => n857);
   U1199 : NAND2X1 port map( A => SUMB_7_5_port, B => n581, Y => n858);
   U1200 : NAND3X1 port map( A => n856, B => n857, C => n858, Y => 
                           CARRYB_8_4_port);
   U1201 : XOR2X1 port map( A => n265, B => ab_14_0_port, Y => n859);
   U1202 : XOR2X1 port map( A => n859, B => n538, Y => A1_12_port);
   U1203 : NAND2X1 port map( A => n546, B => ab_13_1_port, Y => n860);
   U1204 : NAND2X1 port map( A => SUMB_12_2_port, B => ab_13_1_port, Y => n861)
                           ;
   U1205 : NAND2X1 port map( A => SUMB_12_2_port, B => n546, Y => n862);
   U1206 : NAND3X1 port map( A => n860, B => n861, C => n862, Y => 
                           CARRYB_13_1_port);
   U1207 : NAND2X1 port map( A => CARRYB_13_0_port, B => ab_14_0_port, Y => 
                           n863);
   U1208 : NAND2X1 port map( A => SUMB_13_1_port, B => ab_14_0_port, Y => n864)
                           ;
   U1209 : NAND2X1 port map( A => SUMB_13_1_port, B => CARRYB_13_0_port, Y => 
                           n865);
   U1210 : NAND3X1 port map( A => n864, B => n865, C => n863, Y => 
                           CARRYB_14_0_port);
   U1211 : NAND2X1 port map( A => ab_9_7_port, B => n494, Y => n868);
   U1212 : NAND2X1 port map( A => SUMB_8_8_port, B => ab_9_7_port, Y => n869);
   U1213 : NAND2X1 port map( A => SUMB_8_8_port, B => n494, Y => n870);
   U1214 : NAND3X1 port map( A => n868, B => n869, C => n870, Y => 
                           CARRYB_9_7_port);
   U1215 : NAND2X1 port map( A => ab_10_6_port, B => n422, Y => n871);
   U1216 : NAND2X1 port map( A => SUMB_9_7_port, B => ab_10_6_port, Y => n872);
   U1217 : NAND2X1 port map( A => SUMB_9_7_port, B => n422, Y => n873);
   U1218 : NAND3X1 port map( A => n871, B => n872, C => n873, Y => 
                           CARRYB_10_6_port);
   U1219 : XOR2X1 port map( A => n874, B => n43, Y => SUMB_3_13_port);
   U1220 : NAND2X1 port map( A => ab_2_14_port, B => n195, Y => n875);
   U1221 : NAND2X1 port map( A => ab_2_14_port, B => ab_1_15_port, Y => n876);
   U1222 : NAND2X1 port map( A => n195, B => ab_1_15_port, Y => n877);
   U1223 : NAND3X1 port map( A => n875, B => n876, C => n877, Y => 
                           CARRYB_2_14_port);
   U1224 : NAND2X1 port map( A => ab_3_13_port, B => n163, Y => n878);
   U1225 : NAND2X1 port map( A => ab_3_13_port, B => SUMB_2_14_port, Y => n879)
                           ;
   U1226 : NAND2X1 port map( A => n163, B => SUMB_2_14_port, Y => n880);
   U1227 : NAND3X1 port map( A => n878, B => n879, C => n880, Y => 
                           CARRYB_3_13_port);
   U1228 : NAND2X1 port map( A => ab_10_8_port, B => n328, Y => n881);
   U1229 : NAND2X1 port map( A => SUMB_9_9_port, B => ab_10_8_port, Y => n882);
   U1230 : NAND2X1 port map( A => n328, B => SUMB_9_9_port, Y => n883);
   U1231 : NAND3X1 port map( A => n881, B => n882, C => n883, Y => 
                           CARRYB_10_8_port);
   U1232 : NAND2X1 port map( A => ab_11_7_port, B => n658, Y => n884);
   U1233 : NAND2X1 port map( A => SUMB_10_8_port, B => ab_11_7_port, Y => n885)
                           ;
   U1234 : NAND2X1 port map( A => SUMB_10_8_port, B => n658, Y => n886);
   U1235 : NAND3X1 port map( A => n884, B => n885, C => n886, Y => 
                           CARRYB_11_7_port);
   U1236 : XOR2X1 port map( A => ab_13_5_port, B => CARRYB_12_5_port, Y => n887
                           );
   U1237 : XOR2X1 port map( A => n887, B => SUMB_12_6_port, Y => SUMB_13_5_port
                           );
   U1238 : NAND2X1 port map( A => ab_13_5_port, B => CARRYB_12_5_port, Y => 
                           n888);
   U1239 : NAND2X1 port map( A => SUMB_12_6_port, B => ab_13_5_port, Y => n889)
                           ;
   U1240 : NAND2X1 port map( A => SUMB_12_6_port, B => CARRYB_12_5_port, Y => 
                           n890);
   U1241 : NAND3X1 port map( A => n888, B => n889, C => n890, Y => 
                           CARRYB_13_5_port);
   U1242 : NAND2X1 port map( A => ab_14_4_port, B => n495, Y => n891);
   U1243 : NAND2X1 port map( A => SUMB_13_5_port, B => ab_14_4_port, Y => n892)
                           ;
   U1244 : NAND2X1 port map( A => n495, B => SUMB_13_5_port, Y => n893);
   U1245 : NAND3X1 port map( A => n891, B => n892, C => n893, Y => 
                           CARRYB_14_4_port);
   U1246 : INVX1 port map( A => n1061, Y => n894);
   U1247 : NAND2X1 port map( A => ab_9_5_port, B => n393, Y => n895);
   U1248 : NAND2X1 port map( A => SUMB_8_6_port, B => ab_9_5_port, Y => n896);
   U1249 : NAND2X1 port map( A => n393, B => SUMB_8_6_port, Y => n897);
   U1250 : NAND3X1 port map( A => n895, B => n896, C => n897, Y => 
                           CARRYB_9_5_port);
   U1251 : NAND2X1 port map( A => ab_10_4_port, B => n455, Y => n898);
   U1252 : NAND2X1 port map( A => SUMB_9_5_port, B => ab_10_4_port, Y => n899);
   U1253 : NAND2X1 port map( A => SUMB_9_5_port, B => n455, Y => n900);
   U1254 : NAND3X1 port map( A => n898, B => n900, C => n899, Y => 
                           CARRYB_10_4_port);
   U1255 : NAND2X1 port map( A => ab_6_7_port, B => n679, Y => n901);
   U1256 : NAND2X1 port map( A => SUMB_5_8_port, B => ab_6_7_port, Y => n902);
   U1257 : NAND2X1 port map( A => SUMB_5_8_port, B => n679, Y => n903);
   U1258 : NAND3X1 port map( A => n901, B => n903, C => n902, Y => 
                           CARRYB_6_7_port);
   U1259 : NAND2X1 port map( A => ab_7_6_port, B => n125, Y => n904);
   U1260 : NAND2X1 port map( A => SUMB_6_7_port, B => ab_7_6_port, Y => n905);
   U1261 : NAND2X1 port map( A => SUMB_6_7_port, B => n125, Y => n906);
   U1262 : NAND3X1 port map( A => n904, B => n905, C => n906, Y => 
                           CARRYB_7_6_port);
   U1263 : NAND2X1 port map( A => ab_9_4_port, B => n322, Y => n907);
   U1264 : NAND2X1 port map( A => SUMB_8_5_port, B => ab_9_4_port, Y => n908);
   U1265 : NAND2X1 port map( A => SUMB_8_5_port, B => n322, Y => n909);
   U1266 : NAND3X1 port map( A => n907, B => n908, C => n909, Y => 
                           CARRYB_9_4_port);
   U1267 : NAND2X1 port map( A => n317, B => ab_10_3_port, Y => n910);
   U1268 : NAND2X1 port map( A => SUMB_9_4_port, B => ab_10_3_port, Y => n911);
   U1269 : NAND2X1 port map( A => SUMB_9_4_port, B => n317, Y => n912);
   U1270 : NAND3X1 port map( A => n910, B => n911, C => n912, Y => 
                           CARRYB_10_3_port);
   U1271 : INVX2 port map( A => CARRYB_3_8_port, Y => n913);
   U1272 : NAND2X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, Y => n915)
                           ;
   U1273 : NAND2X1 port map( A => SUMB_3_7_port, B => ab_4_6_port, Y => n916);
   U1274 : NAND2X1 port map( A => SUMB_3_7_port, B => CARRYB_3_6_port, Y => 
                           n917);
   U1275 : NAND3X1 port map( A => n915, B => n916, C => n917, Y => 
                           CARRYB_4_6_port);
   U1276 : NAND2X1 port map( A => ab_5_5_port, B => n571, Y => n918);
   U1277 : NAND2X1 port map( A => SUMB_4_6_port, B => ab_5_5_port, Y => n919);
   U1278 : NAND2X1 port map( A => SUMB_4_6_port, B => n571, Y => n920);
   U1279 : NAND3X1 port map( A => n918, B => n920, C => n919, Y => 
                           CARRYB_5_5_port);
   U1280 : NAND2X1 port map( A => SUMB_9_3_port, B => n124, Y => n921);
   U1281 : NAND2X1 port map( A => SUMB_9_3_port, B => ab_10_2_port, Y => n922);
   U1282 : NAND2X1 port map( A => n124, B => ab_10_2_port, Y => n923);
   U1283 : XOR2X1 port map( A => n100, B => n924, Y => SUMB_5_6_port);
   U1284 : NAND2X1 port map( A => ab_4_7_port, B => n655, Y => n925);
   U1285 : NAND2X1 port map( A => SUMB_3_8_port, B => ab_4_7_port, Y => n926);
   U1286 : NAND2X1 port map( A => SUMB_3_8_port, B => n655, Y => n927);
   U1287 : NAND3X1 port map( A => n926, B => n925, C => n927, Y => 
                           CARRYB_4_7_port);
   U1288 : NAND2X1 port map( A => SUMB_4_7_port, B => ab_5_6_port, Y => n929);
   U1289 : NAND2X1 port map( A => SUMB_4_7_port, B => CARRYB_4_6_port, Y => 
                           n930);
   U1290 : NAND3X1 port map( A => n928, B => n929, C => n930, Y => 
                           CARRYB_5_6_port);
   U1291 : NAND2X1 port map( A => SUMB_8_4_port, B => n723, Y => n931);
   U1292 : NAND2X1 port map( A => SUMB_8_4_port, B => ab_9_3_port, Y => n932);
   U1293 : NAND2X1 port map( A => n723, B => ab_9_3_port, Y => n933);
   U1294 : NAND3X1 port map( A => n933, B => n931, C => n932, Y => 
                           CARRYB_9_3_port);
   U1295 : NAND2X1 port map( A => n3, B => ab_2_8_port, Y => n934);
   U1296 : NAND2X1 port map( A => SUMB_1_9_port, B => ab_2_8_port, Y => n935);
   U1297 : NAND2X1 port map( A => SUMB_1_9_port, B => n3, Y => n936);
   U1298 : NAND3X1 port map( A => n934, B => n935, C => n936, Y => 
                           CARRYB_2_8_port);
   U1299 : NAND2X1 port map( A => ab_3_7_port, B => n391, Y => n937);
   U1300 : NAND2X1 port map( A => SUMB_2_8_port, B => ab_3_7_port, Y => n938);
   U1301 : NAND2X1 port map( A => SUMB_2_8_port, B => n391, Y => n939);
   U1302 : NAND3X1 port map( A => n937, B => n938, C => n939, Y => 
                           CARRYB_3_7_port);
   U1303 : NAND2X1 port map( A => ab_6_8_port, B => n946, Y => n940);
   U1304 : NAND2X1 port map( A => SUMB_5_9_port, B => ab_6_8_port, Y => n941);
   U1305 : NAND2X1 port map( A => SUMB_5_9_port, B => n946, Y => n942);
   U1306 : NAND3X1 port map( A => n940, B => n941, C => n942, Y => 
                           CARRYB_6_8_port);
   U1307 : NAND2X1 port map( A => n792, B => ab_7_7_port, Y => n943);
   U1308 : NAND2X1 port map( A => SUMB_6_8_port, B => ab_7_7_port, Y => n944);
   U1309 : NAND2X1 port map( A => SUMB_6_8_port, B => n792, Y => n945);
   U1310 : NAND3X1 port map( A => n944, B => n943, C => n945, Y => 
                           CARRYB_7_7_port);
   U1311 : NAND2X1 port map( A => ab_2_5_port, B => n439, Y => n948);
   U1312 : NAND2X1 port map( A => ab_2_5_port, B => SUMB_1_6_port, Y => n949);
   U1313 : NAND2X1 port map( A => n439, B => SUMB_1_6_port, Y => n950);
   U1314 : NAND3X1 port map( A => n948, B => n949, C => n950, Y => 
                           CARRYB_2_5_port);
   U1315 : NAND2X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, Y => n951)
                           ;
   U1316 : NAND2X1 port map( A => ab_3_4_port, B => SUMB_2_5_port, Y => n952);
   U1317 : NAND2X1 port map( A => CARRYB_2_4_port, B => SUMB_2_5_port, Y => 
                           n953);
   U1318 : NAND3X1 port map( A => n951, B => n952, C => n953, Y => 
                           CARRYB_3_4_port);
   U1319 : XNOR2X1 port map( A => CARRYB_14_0_port, B => ab_15_0_port, Y => 
                           n954);
   U1320 : XOR2X1 port map( A => CARRYB_7_7_port, B => ab_8_7_port, Y => n955);
   U1321 : XOR2X1 port map( A => SUMB_7_8_port, B => n955, Y => SUMB_8_7_port);
   U1322 : NAND2X1 port map( A => ab_8_7_port, B => n969, Y => n957);
   U1323 : NAND2X1 port map( A => SUMB_7_8_port, B => ab_8_7_port, Y => n958);
   U1324 : NAND2X1 port map( A => SUMB_7_8_port, B => n969, Y => n959);
   U1325 : NAND3X1 port map( A => n957, B => n958, C => n959, Y => 
                           CARRYB_8_7_port);
   U1326 : NAND2X1 port map( A => ab_9_6_port, B => n130, Y => n960);
   U1327 : NAND2X1 port map( A => SUMB_8_7_port, B => ab_9_6_port, Y => n961);
   U1328 : NAND2X1 port map( A => n130, B => SUMB_8_7_port, Y => n962);
   U1329 : NAND3X1 port map( A => n960, B => n961, C => n962, Y => 
                           CARRYB_9_6_port);
   U1330 : NAND2X1 port map( A => ab_14_1_port, B => n1031, Y => n963);
   U1331 : NAND2X1 port map( A => SUMB_13_2_port, B => ab_14_1_port, Y => n964)
                           ;
   U1332 : NAND2X1 port map( A => SUMB_13_2_port, B => n1031, Y => n965);
   U1333 : NAND3X1 port map( A => n965, B => n963, C => n964, Y => 
                           CARRYB_14_1_port);
   U1334 : NAND2X1 port map( A => n418, B => ab_15_0_port, Y => n966);
   U1335 : NAND2X1 port map( A => ab_15_0_port, B => SUMB_14_1_port, Y => n967)
                           ;
   U1336 : NAND2X1 port map( A => n418, B => SUMB_14_1_port, Y => n968);
   U1337 : NAND3X1 port map( A => n966, B => n968, C => n967, Y => 
                           CARRYB_15_0_port);
   U1338 : NAND2X1 port map( A => CARRYB_6_4_port, B => ab_7_4_port, Y => n970)
                           ;
   U1339 : NAND2X1 port map( A => SUMB_6_5_port, B => ab_7_4_port, Y => n971);
   U1340 : NAND2X1 port map( A => SUMB_6_5_port, B => n420, Y => n972);
   U1341 : NAND3X1 port map( A => n970, B => n971, C => n972, Y => 
                           CARRYB_7_4_port);
   U1342 : NAND2X1 port map( A => ab_8_3_port, B => n141, Y => n973);
   U1343 : NAND2X1 port map( A => SUMB_7_4_port, B => ab_8_3_port, Y => n974);
   U1344 : NAND2X1 port map( A => n348, B => SUMB_7_4_port, Y => n975);
   U1345 : NAND3X1 port map( A => n18, B => n974, C => n975, Y => 
                           CARRYB_8_3_port);
   U1346 : XOR2X1 port map( A => n210, B => ab_2_6_port, Y => n976);
   U1347 : NAND2X1 port map( A => n210, B => ab_2_6_port, Y => n977);
   U1348 : NAND2X1 port map( A => ab_2_6_port, B => SUMB_1_7_port, Y => n978);
   U1349 : NAND2X1 port map( A => n210, B => SUMB_1_7_port, Y => n979);
   U1350 : NAND3X1 port map( A => n977, B => n978, C => n979, Y => 
                           CARRYB_2_6_port);
   U1351 : NAND2X1 port map( A => ab_3_5_port, B => n986, Y => n980);
   U1352 : NAND2X1 port map( A => SUMB_2_6_port, B => ab_3_5_port, Y => n981);
   U1353 : NAND2X1 port map( A => SUMB_2_6_port, B => n986, Y => n982);
   U1354 : NAND3X1 port map( A => n980, B => n981, C => n982, Y => 
                           CARRYB_3_5_port);
   U1355 : INVX2 port map( A => CARRYB_2_5_port, Y => n985);
   U1356 : XOR2X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, Y => n987);
   U1357 : XOR2X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, Y => n988);
   U1358 : XOR2X1 port map( A => n988, B => n476, Y => SUMB_4_2_port);
   U1359 : NAND2X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, Y => n989)
                           ;
   U1360 : NAND2X1 port map( A => ab_3_3_port, B => SUMB_2_4_port, Y => n990);
   U1361 : NAND2X1 port map( A => CARRYB_2_3_port, B => SUMB_2_4_port, Y => 
                           n991);
   U1362 : NAND3X1 port map( A => n989, B => n990, C => n991, Y => 
                           CARRYB_3_3_port);
   U1363 : NAND2X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, Y => n992)
                           ;
   U1364 : NAND2X1 port map( A => ab_4_2_port, B => SUMB_3_3_port, Y => n993);
   U1365 : NAND2X1 port map( A => CARRYB_3_2_port, B => SUMB_3_3_port, Y => 
                           n994);
   U1366 : NAND3X1 port map( A => n992, B => n993, C => n994, Y => 
                           CARRYB_4_2_port);
   U1367 : XOR2X1 port map( A => n427, B => ab_7_1_port, Y => n995);
   U1368 : XOR2X1 port map( A => n995, B => n1003, Y => SUMB_7_1_port);
   U1369 : XOR2X1 port map( A => ab_8_0_port, B => n140, Y => n996);
   U1370 : XOR2X1 port map( A => n996, B => SUMB_7_1_port, Y => A1_6_port);
   U1371 : NAND2X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, Y => n997)
                           ;
   U1372 : NAND2X1 port map( A => ab_7_1_port, B => SUMB_6_2_port, Y => n998);
   U1373 : NAND2X1 port map( A => SUMB_6_2_port, B => CARRYB_6_1_port, Y => 
                           n999);
   U1374 : NAND3X1 port map( A => n998, B => n997, C => n999, Y => 
                           CARRYB_7_1_port);
   U1375 : NAND2X1 port map( A => ab_8_0_port, B => CARRYB_7_0_port, Y => n1000
                           );
   U1376 : NAND2X1 port map( A => ab_8_0_port, B => SUMB_7_1_port, Y => n1001);
   U1377 : NAND2X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Y => 
                           n1002);
   U1378 : NAND3X1 port map( A => n1002, B => n1001, C => n1000, Y => 
                           CARRYB_8_0_port);
   U1379 : BUFX2 port map( A => SUMB_6_2_port, Y => n1003);
   U1380 : XOR2X1 port map( A => CARRYB_2_2_port, B => ab_3_2_port, Y => n1004)
                           ;
   U1381 : XOR2X1 port map( A => n624, B => n1004, Y => SUMB_3_2_port);
   U1382 : NAND2X1 port map( A => SUMB_2_3_port, B => CARRYB_2_2_port, Y => 
                           n1005);
   U1383 : NAND2X1 port map( A => SUMB_2_3_port, B => ab_3_2_port, Y => n1006);
   U1384 : NAND2X1 port map( A => CARRYB_2_2_port, B => ab_3_2_port, Y => n1007
                           );
   U1385 : NAND3X1 port map( A => n1006, B => n1005, C => n1007, Y => 
                           CARRYB_3_2_port);
   U1386 : NAND2X1 port map( A => SUMB_6_3_port, B => ab_7_2_port, Y => n1009);
   U1387 : NAND2X1 port map( A => n5, B => SUMB_6_3_port, Y => n1010);
   U1388 : NAND3X1 port map( A => n423, B => n1009, C => n1010, Y => 
                           CARRYB_7_2_port);
   U1389 : NAND2X1 port map( A => CARRYB_7_1_port, B => ab_8_1_port, Y => n1011
                           );
   U1390 : NAND2X1 port map( A => SUMB_7_2_port, B => ab_8_1_port, Y => n1012);
   U1391 : NAND2X1 port map( A => SUMB_7_2_port, B => CARRYB_7_1_port, Y => 
                           n1013);
   U1392 : NAND3X1 port map( A => n1011, B => n1012, C => n1013, Y => 
                           CARRYB_8_1_port);
   U1393 : INVX4 port map( A => A(0), Y => n1061);
   U1394 : AND2X2 port map( A => SUMB_15_1_port, B => n115, Y => n1014);
   U1395 : AND2X2 port map( A => SUMB_15_2_port, B => CARRYB_15_1_port, Y => 
                           n1015);
   U1396 : AND2X2 port map( A => ab_0_1_port, B => ab_1_0_port, Y => n1020);
   U1397 : INVX1 port map( A => B(1), Y => n1034);
   U1398 : INVX2 port map( A => B(10), Y => n1051);
   U1399 : INVX2 port map( A => A(13), Y => n1098);
   U1400 : INVX2 port map( A => A(15), Y => n1096);
   U1401 : INVX2 port map( A => A(14), Y => n1097);
   U1402 : INVX2 port map( A => A(4), Y => n1068);
   U1403 : INVX2 port map( A => A(5), Y => n1070);
   U1404 : INVX2 port map( A => A(6), Y => n1072);
   U1405 : INVX2 port map( A => A(7), Y => n1074);
   U1406 : INVX2 port map( A => A(9), Y => n1078);
   U1407 : INVX2 port map( A => A(8), Y => n1076);
   U1408 : INVX2 port map( A => A(10), Y => n1080);
   U1409 : XOR2X1 port map( A => SUMB_15_2_port, B => CARRYB_15_1_port, Y => 
                           A1_15_port);
   U1410 : XOR2X1 port map( A => SUMB_15_3_port, B => CARRYB_15_2_port, Y => 
                           A1_16_port);
   U1411 : XOR2X1 port map( A => SUMB_15_4_port, B => CARRYB_15_3_port, Y => 
                           A1_17_port);
   U1412 : XOR2X1 port map( A => SUMB_15_5_port, B => CARRYB_15_4_port, Y => 
                           A1_18_port);
   U1413 : NAND2X1 port map( A => SUMB_15_7_port, B => CARRYB_15_6_port, Y => 
                           n1023);
   U1414 : INVX2 port map( A => n1023, Y => A2_21_port);
   U1415 : XOR2X1 port map( A => SUMB_15_8_port, B => CARRYB_15_7_port, Y => 
                           A1_21_port);
   U1416 : XOR2X1 port map( A => SUMB_15_9_port, B => CARRYB_15_8_port, Y => 
                           A1_22_port);
   U1417 : XOR2X1 port map( A => SUMB_15_10_port, B => CARRYB_15_9_port, Y => 
                           A1_23_port);
   U1418 : XOR2X1 port map( A => SUMB_15_11_port, B => CARRYB_15_10_port, Y => 
                           A1_24_port);
   U1419 : XOR2X1 port map( A => SUMB_15_12_port, B => CARRYB_15_11_port, Y => 
                           A1_25_port);
   U1420 : XOR2X1 port map( A => SUMB_15_13_port, B => CARRYB_15_12_port, Y => 
                           A1_26_port);
   U1421 : XOR2X1 port map( A => SUMB_15_14_port, B => CARRYB_15_13_port, Y => 
                           A1_27_port);
   U1422 : XOR2X1 port map( A => SUMB_15_15_port, B => CARRYB_15_14_port, Y => 
                           A1_28_port);
   U1423 : XOR2X1 port map( A => ab_1_0_port, B => ab_0_1_port, Y => PRODUCT(1)
                           );
   U1424 : XOR2X1 port map( A => ab_1_1_port, B => ab_0_2_port, Y => 
                           SUMB_1_1_port);
   U1425 : XOR2X1 port map( A => n1022, B => ab_0_3_port, Y => SUMB_1_2_port);
   U1426 : XOR2X1 port map( A => ab_1_3_port, B => ab_0_4_port, Y => 
                           SUMB_1_3_port);
   U1427 : XOR2X1 port map( A => ab_1_5_port, B => ab_0_6_port, Y => 
                           SUMB_1_5_port);
   U1428 : XOR2X1 port map( A => ab_1_6_port, B => ab_0_7_port, Y => 
                           SUMB_1_6_port);
   U1429 : XOR2X1 port map( A => ab_0_11_port, B => ab_1_10_port, Y => 
                           SUMB_1_10_port);
   U1430 : NAND2X1 port map( A => ab_0_11_port, B => ab_1_10_port, Y => n1024);
   U1431 : XOR2X1 port map( A => ab_1_11_port, B => ab_0_12_port, Y => 
                           SUMB_1_11_port);
   U1432 : XOR2X1 port map( A => ab_0_13_port, B => ab_1_12_port, Y => 
                           SUMB_1_12_port);
   U1433 : XOR2X1 port map( A => ab_1_13_port, B => ab_0_14_port, Y => 
                           SUMB_1_13_port);
   U1434 : NAND2X1 port map( A => ab_0_14_port, B => ab_1_13_port, Y => n1025);
   U1435 : INVX2 port map( A => n1025, Y => CARRYB_1_13_port);
   U1436 : XOR2X1 port map( A => ab_1_14_port, B => ab_0_15_port, Y => 
                           SUMB_1_14_port);
   U1437 : BUFX4 port map( A => CARRYB_9_1_port, Y => n1026);
   U1438 : INVX1 port map( A => n1039, Y => n1091);
   U1439 : INVX1 port map( A => n1035, Y => n1093);
   U1440 : INVX2 port map( A => CARRYB_6_2_port, Y => n1027);
   U1441 : INVX1 port map( A => n1041, Y => n1090);
   U1442 : INVX4 port map( A => B(4), Y => n1040);
   U1443 : INVX2 port map( A => CARRYB_10_3_port, Y => n1028);
   U1444 : INVX4 port map( A => B(2), Y => n1036);
   U1445 : INVX2 port map( A => CARRYB_13_1_port, Y => n1030);
   U1446 : INVX8 port map( A => n1032, Y => n1033);
   U1447 : INVX8 port map( A => n1036, Y => n1037);
   U1448 : INVX8 port map( A => n1038, Y => n1039);
   U1449 : INVX8 port map( A => n1040, Y => n1041);
   U1450 : INVX8 port map( A => n1042, Y => n1043);
   U1451 : INVX8 port map( A => n1044, Y => n1045);
   U1452 : INVX8 port map( A => n1051, Y => n1052);
   U1453 : INVX8 port map( A => n1055, Y => n1056);
   U1454 : INVX8 port map( A => n1057, Y => n1058);
   U1455 : INVX8 port map( A => n1059, Y => n1060);
   U1456 : INVX8 port map( A => n1064, Y => n1065);
   U1457 : INVX8 port map( A => n1066, Y => n1067);
   U1458 : INVX8 port map( A => n1068, Y => n1069);
   U1459 : INVX8 port map( A => n1070, Y => n1071);
   U1460 : INVX8 port map( A => n1072, Y => n1073);
   U1461 : INVX8 port map( A => n1074, Y => n1075);
   U1462 : INVX8 port map( A => n1076, Y => n1077);
   U1463 : INVX8 port map( A => n1078, Y => n1079);
   U1464 : AND2X2 port map( A => n42, B => n1060, Y => ab_1_14_port);
   U1465 : AND2X2 port map( A => n1060, B => n103, Y => ab_0_14_port);
   U1466 : AND2X2 port map( A => n983, B => n1058, Y => ab_1_13_port);
   U1467 : AND2X2 port map( A => n1058, B => n1062, Y => ab_0_13_port);
   U1468 : AND2X2 port map( A => n42, B => n1056, Y => ab_1_12_port);
   U1469 : AND2X2 port map( A => n1056, B => n298, Y => ab_0_12_port);
   U1470 : AND2X2 port map( A => n42, B => B(11), Y => ab_1_11_port);
   U1471 : AND2X2 port map( A => n1062, B => B(11), Y => ab_0_11_port);
   U1472 : AND2X2 port map( A => n983, B => n1052, Y => ab_1_10_port);
   U1473 : AND2X2 port map( A => n1052, B => n298, Y => ab_0_10_port);
   U1474 : AND2X2 port map( A => B(7), B => n1062, Y => ab_0_7_port);
   U1475 : AND2X2 port map( A => n983, B => n1043, Y => ab_1_5_port);
   U1476 : AND2X2 port map( A => n1043, B => n103, Y => ab_0_5_port);
   U1477 : AND2X2 port map( A => n1041, B => n983, Y => ab_1_4_port);
   U1478 : AND2X2 port map( A => n1041, B => n103, Y => ab_0_4_port);
   U1479 : AND2X2 port map( A => n1039, B => n984, Y => ab_1_3_port);
   U1480 : AND2X2 port map( A => n1039, B => n105, Y => ab_0_3_port);
   U1481 : AND2X2 port map( A => n1037, B => n894, Y => ab_0_2_port);
   U1482 : AND2X2 port map( A => B(1), B => n894, Y => ab_0_1_port);
   U1483 : AND2X2 port map( A => n984, B => B(0), Y => ab_1_0_port);
   U1484 : AND2X2 port map( A => n1065, B => n1060, Y => ab_2_14_port);
   U1485 : NOR2X1 port map( A => n984, B => n1095, Y => ab_1_15_port);
   U1486 : AND2X2 port map( A => n1065, B => n1058, Y => ab_2_13_port);
   U1487 : AND2X2 port map( A => n1065, B => n1056, Y => ab_2_12_port);
   U1488 : AND2X2 port map( A => n1065, B => B(11), Y => ab_2_11_port);
   U1489 : AND2X2 port map( A => n1065, B => n1052, Y => ab_2_10_port);
   U1490 : AND2X2 port map( A => n1065, B => n579, Y => ab_2_9_port);
   U1491 : AND2X2 port map( A => n1065, B => n529, Y => ab_2_8_port);
   U1492 : AND2X2 port map( A => n1065, B => B(7), Y => ab_2_7_port);
   U1493 : AND2X2 port map( A => n1065, B => n1045, Y => ab_2_6_port);
   U1494 : AND2X2 port map( A => n1065, B => n1043, Y => ab_2_5_port);
   U1495 : AND2X2 port map( A => n1065, B => n1041, Y => ab_2_4_port);
   U1496 : AND2X2 port map( A => n1065, B => n1039, Y => ab_2_3_port);
   U1497 : AND2X2 port map( A => n1065, B => n1037, Y => ab_2_2_port);
   U1498 : AND2X2 port map( A => n153, B => B(1), Y => ab_2_1_port);
   U1499 : AND2X2 port map( A => n153, B => n1033, Y => ab_2_0_port);
   U1500 : AND2X2 port map( A => n1067, B => n1060, Y => ab_3_14_port);
   U1501 : NOR2X1 port map( A => n153, B => n1095, Y => ab_2_15_port);
   U1502 : AND2X2 port map( A => n1067, B => n1058, Y => ab_3_13_port);
   U1503 : AND2X2 port map( A => n1067, B => n1056, Y => ab_3_12_port);
   U1504 : AND2X2 port map( A => n1067, B => B(11), Y => ab_3_11_port);
   U1505 : AND2X2 port map( A => n1067, B => n1052, Y => ab_3_10_port);
   U1506 : AND2X2 port map( A => n1067, B => n579, Y => ab_3_9_port);
   U1507 : AND2X2 port map( A => n1067, B => n529, Y => ab_3_8_port);
   U1508 : AND2X2 port map( A => n1067, B => n1047, Y => ab_3_7_port);
   U1509 : AND2X2 port map( A => n1067, B => n1045, Y => ab_3_6_port);
   U1510 : AND2X2 port map( A => n1067, B => n1043, Y => ab_3_5_port);
   U1511 : AND2X2 port map( A => n1067, B => n1041, Y => ab_3_4_port);
   U1512 : AND2X2 port map( A => n1067, B => n1039, Y => ab_3_3_port);
   U1513 : AND2X2 port map( A => n1067, B => n1037, Y => ab_3_2_port);
   U1514 : AND2X2 port map( A => n1067, B => B(1), Y => ab_3_1_port);
   U1515 : AND2X2 port map( A => n1067, B => n1033, Y => ab_3_0_port);
   U1516 : AND2X2 port map( A => n1069, B => n1060, Y => ab_4_14_port);
   U1517 : NOR2X1 port map( A => n1067, B => n1095, Y => ab_3_15_port);
   U1518 : AND2X2 port map( A => n1069, B => n1058, Y => ab_4_13_port);
   U1519 : AND2X2 port map( A => n1069, B => n1056, Y => ab_4_12_port);
   U1520 : AND2X2 port map( A => n1069, B => n1054, Y => ab_4_11_port);
   U1521 : AND2X2 port map( A => n1069, B => n1052, Y => ab_4_10_port);
   U1522 : AND2X2 port map( A => n1069, B => n579, Y => ab_4_9_port);
   U1523 : AND2X2 port map( A => n1069, B => n529, Y => ab_4_8_port);
   U1524 : AND2X2 port map( A => n1069, B => n1047, Y => ab_4_7_port);
   U1525 : AND2X2 port map( A => n1069, B => n1045, Y => ab_4_6_port);
   U1526 : AND2X2 port map( A => n1069, B => n1043, Y => ab_4_5_port);
   U1527 : AND2X2 port map( A => n1069, B => n1041, Y => ab_4_4_port);
   U1528 : AND2X2 port map( A => n1069, B => n1039, Y => ab_4_3_port);
   U1529 : AND2X2 port map( A => n1069, B => n1037, Y => ab_4_2_port);
   U1530 : AND2X2 port map( A => n1069, B => n1035, Y => ab_4_1_port);
   U1531 : AND2X2 port map( A => n1069, B => n1033, Y => ab_4_0_port);
   U1532 : AND2X2 port map( A => n1071, B => n1060, Y => ab_5_14_port);
   U1533 : NOR2X1 port map( A => n1069, B => n1095, Y => ab_4_15_port);
   U1534 : AND2X2 port map( A => n1071, B => n1058, Y => ab_5_13_port);
   U1535 : AND2X2 port map( A => n1071, B => n1056, Y => ab_5_12_port);
   U1536 : AND2X2 port map( A => n1071, B => n1054, Y => ab_5_11_port);
   U1537 : AND2X2 port map( A => n1071, B => n1052, Y => ab_5_10_port);
   U1538 : AND2X2 port map( A => n1071, B => n579, Y => ab_5_9_port);
   U1539 : AND2X2 port map( A => n1071, B => n529, Y => ab_5_8_port);
   U1540 : AND2X2 port map( A => n1071, B => n1047, Y => ab_5_7_port);
   U1541 : AND2X2 port map( A => n1071, B => n1045, Y => ab_5_6_port);
   U1542 : AND2X2 port map( A => n1071, B => n1043, Y => ab_5_5_port);
   U1543 : AND2X2 port map( A => n1071, B => n1041, Y => ab_5_4_port);
   U1544 : AND2X2 port map( A => n1071, B => n1039, Y => ab_5_3_port);
   U1545 : AND2X2 port map( A => n1071, B => n1037, Y => ab_5_2_port);
   U1546 : AND2X2 port map( A => n1071, B => n1035, Y => ab_5_1_port);
   U1547 : AND2X2 port map( A => n1071, B => n1033, Y => ab_5_0_port);
   U1548 : AND2X2 port map( A => n1073, B => n1060, Y => ab_6_14_port);
   U1549 : NOR2X1 port map( A => n1071, B => n1095, Y => ab_5_15_port);
   U1550 : AND2X2 port map( A => n1073, B => n1058, Y => ab_6_13_port);
   U1551 : AND2X2 port map( A => n1073, B => n1056, Y => ab_6_12_port);
   U1552 : AND2X2 port map( A => n1073, B => n1054, Y => ab_6_11_port);
   U1553 : AND2X2 port map( A => n1073, B => n1052, Y => ab_6_10_port);
   U1554 : AND2X2 port map( A => n1073, B => n579, Y => ab_6_9_port);
   U1555 : AND2X2 port map( A => n1073, B => n529, Y => ab_6_8_port);
   U1556 : AND2X2 port map( A => n1073, B => n1047, Y => ab_6_7_port);
   U1557 : AND2X2 port map( A => n1073, B => n1045, Y => ab_6_6_port);
   U1558 : AND2X2 port map( A => n1073, B => n1043, Y => ab_6_5_port);
   U1559 : AND2X2 port map( A => n1073, B => n1041, Y => ab_6_4_port);
   U1560 : AND2X2 port map( A => n1073, B => n1039, Y => ab_6_3_port);
   U1561 : AND2X2 port map( A => n1073, B => n1037, Y => ab_6_2_port);
   U1562 : AND2X2 port map( A => n1073, B => n1035, Y => ab_6_1_port);
   U1563 : AND2X2 port map( A => n1073, B => n1033, Y => ab_6_0_port);
   U1564 : AND2X2 port map( A => n1075, B => n1060, Y => ab_7_14_port);
   U1565 : NOR2X1 port map( A => n1073, B => n1095, Y => ab_6_15_port);
   U1566 : AND2X2 port map( A => n1075, B => n1058, Y => ab_7_13_port);
   U1567 : AND2X2 port map( A => n1075, B => n1056, Y => ab_7_12_port);
   U1568 : AND2X2 port map( A => n1075, B => n1054, Y => ab_7_11_port);
   U1569 : AND2X2 port map( A => n1075, B => n1052, Y => ab_7_10_port);
   U1570 : AND2X2 port map( A => n1075, B => n579, Y => ab_7_9_port);
   U1571 : AND2X2 port map( A => n1075, B => n529, Y => ab_7_8_port);
   U1572 : AND2X2 port map( A => n1075, B => n1047, Y => ab_7_7_port);
   U1573 : AND2X2 port map( A => n1075, B => n1045, Y => ab_7_6_port);
   U1574 : AND2X2 port map( A => n1075, B => n1043, Y => ab_7_5_port);
   U1575 : AND2X2 port map( A => n1075, B => n1041, Y => ab_7_4_port);
   U1576 : AND2X2 port map( A => n1075, B => n1039, Y => ab_7_3_port);
   U1577 : AND2X2 port map( A => n1075, B => n1037, Y => ab_7_2_port);
   U1578 : AND2X2 port map( A => n1075, B => n1035, Y => ab_7_1_port);
   U1579 : AND2X2 port map( A => n1075, B => n1033, Y => ab_7_0_port);
   U1580 : AND2X2 port map( A => n1077, B => n1060, Y => ab_8_14_port);
   U1581 : NOR2X1 port map( A => n1075, B => n1095, Y => ab_7_15_port);
   U1582 : AND2X2 port map( A => n1077, B => n1058, Y => ab_8_13_port);
   U1583 : AND2X2 port map( A => n1077, B => n1056, Y => ab_8_12_port);
   U1584 : AND2X2 port map( A => n1077, B => n1054, Y => ab_8_11_port);
   U1585 : AND2X2 port map( A => n1077, B => n1052, Y => ab_8_10_port);
   U1586 : AND2X2 port map( A => n1077, B => n579, Y => ab_8_9_port);
   U1587 : AND2X2 port map( A => n1077, B => n529, Y => ab_8_8_port);
   U1588 : AND2X2 port map( A => n1077, B => n1047, Y => ab_8_7_port);
   U1589 : AND2X2 port map( A => n1077, B => n1045, Y => ab_8_6_port);
   U1590 : AND2X2 port map( A => n1077, B => n1043, Y => ab_8_5_port);
   U1591 : AND2X2 port map( A => n1077, B => n1041, Y => ab_8_4_port);
   U1592 : AND2X2 port map( A => n1077, B => n1039, Y => ab_8_3_port);
   U1593 : AND2X2 port map( A => n1077, B => n1037, Y => ab_8_2_port);
   U1594 : AND2X2 port map( A => n1077, B => n1035, Y => ab_8_1_port);
   U1595 : AND2X2 port map( A => n1077, B => n1033, Y => ab_8_0_port);
   U1596 : AND2X2 port map( A => n1079, B => n1060, Y => ab_9_14_port);
   U1597 : NOR2X1 port map( A => n1077, B => n1095, Y => ab_8_15_port);
   U1598 : AND2X2 port map( A => n1079, B => n1058, Y => ab_9_13_port);
   U1599 : AND2X2 port map( A => n1079, B => n1056, Y => ab_9_12_port);
   U1600 : AND2X2 port map( A => n1079, B => n1054, Y => ab_9_11_port);
   U1601 : AND2X2 port map( A => n1079, B => n1052, Y => ab_9_10_port);
   U1602 : AND2X2 port map( A => n1079, B => n579, Y => ab_9_9_port);
   U1603 : AND2X2 port map( A => n1079, B => n529, Y => ab_9_8_port);
   U1604 : AND2X2 port map( A => n1079, B => n1047, Y => ab_9_7_port);
   U1605 : AND2X2 port map( A => n1079, B => n1045, Y => ab_9_6_port);
   U1606 : AND2X2 port map( A => n1079, B => n1043, Y => ab_9_5_port);
   U1607 : AND2X2 port map( A => n1079, B => n1041, Y => ab_9_4_port);
   U1608 : AND2X2 port map( A => n1079, B => n1039, Y => ab_9_3_port);
   U1609 : AND2X2 port map( A => n1079, B => n1037, Y => ab_9_2_port);
   U1610 : AND2X2 port map( A => n1079, B => n1035, Y => ab_9_1_port);
   U1611 : AND2X2 port map( A => n1079, B => n1033, Y => ab_9_0_port);
   U1612 : AND2X2 port map( A => n1081, B => n1060, Y => ab_10_14_port);
   U1613 : NOR2X1 port map( A => n1079, B => n1095, Y => ab_9_15_port);
   U1614 : AND2X2 port map( A => n1081, B => n1058, Y => ab_10_13_port);
   U1615 : AND2X2 port map( A => n1081, B => n1056, Y => ab_10_12_port);
   U1616 : AND2X2 port map( A => n1081, B => n1054, Y => ab_10_11_port);
   U1617 : AND2X2 port map( A => n1081, B => n1052, Y => ab_10_10_port);
   U1618 : AND2X2 port map( A => n1081, B => n579, Y => ab_10_9_port);
   U1619 : AND2X2 port map( A => n1081, B => n529, Y => ab_10_8_port);
   U1620 : AND2X2 port map( A => n1081, B => n1047, Y => ab_10_7_port);
   U1621 : AND2X2 port map( A => n1081, B => n1045, Y => ab_10_6_port);
   U1622 : AND2X2 port map( A => n1081, B => n1043, Y => ab_10_5_port);
   U1623 : AND2X2 port map( A => n1081, B => n1041, Y => ab_10_4_port);
   U1624 : AND2X2 port map( A => n1081, B => n1039, Y => ab_10_3_port);
   U1625 : AND2X2 port map( A => n1081, B => n1037, Y => ab_10_2_port);
   U1626 : AND2X2 port map( A => n1081, B => n1035, Y => ab_10_1_port);
   U1627 : AND2X2 port map( A => n1081, B => n1033, Y => ab_10_0_port);
   U1628 : AND2X2 port map( A => A(11), B => n1060, Y => ab_11_14_port);
   U1629 : NOR2X1 port map( A => n1081, B => n1095, Y => ab_10_15_port);
   U1630 : AND2X2 port map( A => A(11), B => n1058, Y => ab_11_13_port);
   U1631 : AND2X2 port map( A => A(11), B => n1056, Y => ab_11_12_port);
   U1632 : AND2X2 port map( A => A(11), B => n1054, Y => ab_11_11_port);
   U1633 : AND2X2 port map( A => A(11), B => n1052, Y => ab_11_10_port);
   U1634 : AND2X2 port map( A => A(11), B => n579, Y => ab_11_9_port);
   U1635 : AND2X2 port map( A => A(11), B => n529, Y => ab_11_8_port);
   U1636 : AND2X2 port map( A => A(11), B => n1047, Y => ab_11_7_port);
   U1637 : AND2X2 port map( A => A(11), B => n1045, Y => ab_11_6_port);
   U1638 : AND2X2 port map( A => A(11), B => n1043, Y => ab_11_5_port);
   U1639 : AND2X2 port map( A => A(11), B => n1041, Y => ab_11_4_port);
   U1640 : AND2X2 port map( A => A(11), B => n1039, Y => ab_11_3_port);
   U1641 : AND2X2 port map( A => A(11), B => n1037, Y => ab_11_2_port);
   U1642 : AND2X2 port map( A => A(11), B => n1035, Y => ab_11_1_port);
   U1643 : AND2X2 port map( A => A(11), B => n1033, Y => ab_11_0_port);
   U1644 : AND2X2 port map( A => A(12), B => n1060, Y => ab_12_14_port);
   U1645 : NOR2X1 port map( A => A(11), B => n1095, Y => ab_11_15_port);
   U1646 : AND2X2 port map( A => A(12), B => n1058, Y => ab_12_13_port);
   U1647 : AND2X2 port map( A => A(12), B => n1056, Y => ab_12_12_port);
   U1648 : AND2X2 port map( A => A(12), B => n1054, Y => ab_12_11_port);
   U1649 : AND2X2 port map( A => A(12), B => n1052, Y => ab_12_10_port);
   U1650 : AND2X2 port map( A => A(12), B => n579, Y => ab_12_9_port);
   U1651 : AND2X2 port map( A => A(12), B => n529, Y => ab_12_8_port);
   U1652 : AND2X2 port map( A => A(12), B => n1047, Y => ab_12_7_port);
   U1653 : AND2X2 port map( A => A(12), B => n1045, Y => ab_12_6_port);
   U1654 : AND2X2 port map( A => A(12), B => n1043, Y => ab_12_5_port);
   U1655 : AND2X2 port map( A => A(12), B => n1041, Y => ab_12_4_port);
   U1656 : AND2X2 port map( A => A(12), B => n1039, Y => ab_12_3_port);
   U1657 : AND2X2 port map( A => A(12), B => n1037, Y => ab_12_2_port);
   U1658 : AND2X2 port map( A => A(12), B => n1035, Y => ab_12_1_port);
   U1659 : AND2X2 port map( A => A(12), B => n1033, Y => ab_12_0_port);
   U1660 : NOR2X1 port map( A => n1098, B => n1082, Y => ab_13_14_port);
   U1661 : NOR2X1 port map( A => A(12), B => n1095, Y => ab_12_15_port);
   U1662 : INVX2 port map( A => n1058, Y => n1083);
   U1663 : NOR2X1 port map( A => n1098, B => n1083, Y => ab_13_13_port);
   U1664 : NOR2X1 port map( A => n1098, B => n1084, Y => ab_13_12_port);
   U1665 : NOR2X1 port map( A => n1098, B => n1053, Y => ab_13_11_port);
   U1666 : NOR2X1 port map( A => n1098, B => n1085, Y => ab_13_10_port);
   U1667 : NOR2X1 port map( A => n1098, B => n1086, Y => ab_13_9_port);
   U1668 : NOR2X1 port map( A => n1098, B => n1048, Y => ab_13_8_port);
   U1669 : NOR2X1 port map( A => n1098, B => n1087, Y => ab_13_7_port);
   U1670 : NOR2X1 port map( A => n1098, B => n1088, Y => ab_13_6_port);
   U1671 : NOR2X1 port map( A => n1098, B => n1089, Y => ab_13_5_port);
   U1672 : NOR2X1 port map( A => n1098, B => n1090, Y => ab_13_4_port);
   U1673 : NOR2X1 port map( A => n1098, B => n1091, Y => ab_13_3_port);
   U1674 : NOR2X1 port map( A => n1098, B => n1092, Y => ab_13_2_port);
   U1675 : NOR2X1 port map( A => n1098, B => n1093, Y => ab_13_1_port);
   U1676 : NOR2X1 port map( A => n1098, B => n1032, Y => ab_13_0_port);
   U1677 : NOR2X1 port map( A => n1097, B => n1082, Y => ab_14_14_port);
   U1678 : NOR2X1 port map( A => A(13), B => n1095, Y => ab_13_15_port);
   U1679 : NOR2X1 port map( A => n1097, B => n1083, Y => ab_14_13_port);
   U1680 : NOR2X1 port map( A => n1097, B => n1084, Y => ab_14_12_port);
   U1681 : NOR2X1 port map( A => n1097, B => n1053, Y => ab_14_11_port);
   U1682 : NOR2X1 port map( A => n1097, B => n1085, Y => ab_14_10_port);
   U1683 : NOR2X1 port map( A => n1097, B => n1086, Y => ab_14_9_port);
   U1684 : NOR2X1 port map( A => n1097, B => n1048, Y => ab_14_8_port);
   U1685 : NOR2X1 port map( A => n1097, B => n1087, Y => ab_14_7_port);
   U1686 : NOR2X1 port map( A => n1097, B => n1088, Y => ab_14_6_port);
   U1687 : NOR2X1 port map( A => n1097, B => n1089, Y => ab_14_5_port);
   U1688 : NOR2X1 port map( A => n1097, B => n1090, Y => ab_14_4_port);
   U1689 : NOR2X1 port map( A => n1097, B => n1091, Y => ab_14_3_port);
   U1690 : NOR2X1 port map( A => n1097, B => n1092, Y => ab_14_2_port);
   U1691 : NOR2X1 port map( A => n1097, B => n1093, Y => ab_14_1_port);
   U1692 : NOR2X1 port map( A => n1097, B => n1032, Y => ab_14_0_port);
   U1693 : NOR2X1 port map( A => n1096, B => n1095, Y => ab_15_15_port);
   U1694 : NOR2X1 port map( A => A(14), B => n1095, Y => ab_14_15_port);
   U1695 : AND2X2 port map( A => n1033, B => n894, Y => PRODUCT(0));
   U1696 : INVX2 port map( A => CARRYB_15_15_port, Y => n1094);
   U1697 : NOR2X1 port map( A => n579, B => n1096, Y => ab_15_9_port);
   U1698 : NOR2X1 port map( A => n529, B => n1096, Y => ab_15_8_port);
   U1699 : NOR2X1 port map( A => n1047, B => n1096, Y => ab_15_7_port);
   U1700 : NOR2X1 port map( A => n1045, B => n1096, Y => ab_15_6_port);
   U1701 : NOR2X1 port map( A => n1043, B => n1096, Y => ab_15_5_port);
   U1702 : NOR2X1 port map( A => n1041, B => n1096, Y => ab_15_4_port);
   U1703 : NOR2X1 port map( A => n1039, B => n1096, Y => ab_15_3_port);
   U1704 : NOR2X1 port map( A => n1037, B => n1096, Y => ab_15_2_port);
   U1705 : NOR2X1 port map( A => n1035, B => n1096, Y => ab_15_1_port);
   U1706 : NOR2X1 port map( A => n1060, B => n1096, Y => ab_15_14_port);
   U1707 : NOR2X1 port map( A => n1058, B => n1096, Y => ab_15_13_port);
   U1708 : NOR2X1 port map( A => n1056, B => n1096, Y => ab_15_12_port);
   U1709 : NOR2X1 port map( A => n1054, B => n1096, Y => ab_15_11_port);
   U1710 : NOR2X1 port map( A => n1052, B => n1096, Y => ab_15_10_port);
   U1711 : NOR2X1 port map( A => n1033, B => n1096, Y => ab_15_0_port);
   n1099 <= '0';

end SYN_csa;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math_DW02_mult_0 is

   port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  PRODUCT
         : out std_logic_vector (31 downto 0));

end matrix_math_DW02_mult_0;

architecture SYN_csa of matrix_math_DW02_mult_0 is

   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component matrix_math_DW01_add_24
      port( A, B : in std_logic_vector (29 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (29 downto 0);  CO : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_15_15_port, ab_15_14_port, ab_15_13_port, 
      ab_15_12_port, ab_15_11_port, ab_15_10_port, ab_15_9_port, ab_15_8_port, 
      ab_15_7_port, ab_15_6_port, ab_15_5_port, ab_15_4_port, ab_15_3_port, 
      ab_15_2_port, ab_15_1_port, ab_15_0_port, ab_14_15_port, ab_14_14_port, 
      ab_14_13_port, ab_14_12_port, ab_14_11_port, ab_14_10_port, ab_14_9_port,
      ab_14_8_port, ab_14_7_port, ab_14_6_port, ab_14_5_port, ab_14_4_port, 
      ab_14_3_port, ab_14_2_port, ab_14_1_port, ab_14_0_port, ab_13_15_port, 
      ab_13_14_port, ab_13_13_port, ab_13_12_port, ab_13_11_port, ab_13_10_port
      , ab_13_9_port, ab_13_8_port, ab_13_7_port, ab_13_6_port, ab_13_5_port, 
      ab_13_4_port, ab_13_3_port, ab_13_2_port, ab_13_1_port, ab_13_0_port, 
      ab_12_15_port, ab_12_14_port, ab_12_13_port, ab_12_12_port, ab_12_11_port
      , ab_12_10_port, ab_12_9_port, ab_12_8_port, ab_12_7_port, ab_12_6_port, 
      ab_12_5_port, ab_12_4_port, ab_12_3_port, ab_12_2_port, ab_12_1_port, 
      ab_12_0_port, ab_11_15_port, ab_11_14_port, ab_11_13_port, ab_11_12_port,
      ab_11_11_port, ab_11_10_port, ab_11_9_port, ab_11_8_port, ab_11_7_port, 
      ab_11_6_port, ab_11_5_port, ab_11_4_port, ab_11_3_port, ab_11_2_port, 
      ab_11_1_port, ab_11_0_port, ab_10_15_port, ab_10_14_port, ab_10_13_port, 
      ab_10_12_port, ab_10_11_port, ab_10_10_port, ab_10_9_port, ab_10_8_port, 
      ab_10_7_port, ab_10_6_port, ab_10_5_port, ab_10_4_port, ab_10_3_port, 
      ab_10_2_port, ab_10_1_port, ab_10_0_port, ab_9_15_port, ab_9_14_port, 
      ab_9_13_port, ab_9_12_port, ab_9_11_port, ab_9_10_port, ab_9_9_port, 
      ab_9_8_port, ab_9_7_port, ab_9_6_port, ab_9_5_port, ab_9_4_port, 
      ab_9_3_port, ab_9_2_port, ab_9_1_port, ab_9_0_port, ab_8_15_port, 
      ab_8_14_port, ab_8_13_port, ab_8_12_port, ab_8_11_port, ab_8_10_port, 
      ab_8_9_port, ab_8_8_port, ab_8_7_port, ab_8_6_port, ab_8_5_port, 
      ab_8_4_port, ab_8_3_port, ab_8_2_port, ab_8_1_port, ab_8_0_port, 
      ab_7_15_port, ab_7_14_port, ab_7_13_port, ab_7_12_port, ab_7_11_port, 
      ab_7_10_port, ab_7_9_port, ab_7_8_port, ab_7_7_port, ab_7_6_port, 
      ab_7_5_port, ab_7_4_port, ab_7_3_port, ab_7_2_port, ab_7_1_port, 
      ab_7_0_port, ab_6_15_port, ab_6_14_port, ab_6_13_port, ab_6_12_port, 
      ab_6_11_port, ab_6_10_port, ab_6_9_port, ab_6_8_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_15_port, ab_5_14_port, ab_5_13_port, 
      ab_5_12_port, ab_5_11_port, ab_5_10_port, ab_5_9_port, ab_5_8_port, 
      ab_5_7_port, ab_5_6_port, ab_5_5_port, ab_5_4_port, ab_5_3_port, 
      ab_5_2_port, ab_5_1_port, ab_5_0_port, ab_4_15_port, ab_4_14_port, 
      ab_4_13_port, ab_4_12_port, ab_4_11_port, ab_4_10_port, ab_4_9_port, 
      ab_4_8_port, ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, 
      ab_4_3_port, ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_15_port, 
      ab_3_14_port, ab_3_13_port, ab_3_12_port, ab_3_11_port, ab_3_10_port, 
      ab_3_9_port, ab_3_8_port, ab_3_7_port, ab_3_6_port, ab_3_5_port, 
      ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, ab_3_0_port, 
      ab_2_15_port, ab_2_14_port, ab_2_13_port, ab_2_12_port, ab_2_11_port, 
      ab_2_10_port, ab_2_9_port, ab_2_6_port, ab_2_4_port, ab_2_3_port, 
      ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_15_port, ab_1_14_port, 
      ab_1_13_port, ab_1_12_port, ab_1_11_port, ab_1_10_port, ab_1_8_port, 
      ab_1_6_port, ab_1_5_port, ab_1_3_port, ab_1_1_port, ab_1_0_port, 
      ab_0_15_port, ab_0_14_port, ab_0_13_port, ab_0_11_port, ab_0_10_port, 
      ab_0_9_port, ab_0_8_port, ab_0_7_port, ab_0_5_port, ab_0_4_port, 
      ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_15_15_port, 
      CARRYB_15_14_port, CARRYB_15_13_port, CARRYB_15_12_port, 
      CARRYB_15_11_port, CARRYB_15_10_port, CARRYB_15_9_port, CARRYB_15_8_port,
      CARRYB_15_7_port, CARRYB_15_6_port, CARRYB_15_5_port, CARRYB_15_4_port, 
      CARRYB_15_3_port, CARRYB_15_2_port, CARRYB_15_1_port, CARRYB_15_0_port, 
      CARRYB_14_14_port, CARRYB_14_13_port, CARRYB_14_12_port, 
      CARRYB_14_11_port, CARRYB_14_10_port, CARRYB_14_9_port, CARRYB_14_8_port,
      CARRYB_14_7_port, CARRYB_14_6_port, CARRYB_14_5_port, CARRYB_14_4_port, 
      CARRYB_14_3_port, CARRYB_14_2_port, CARRYB_14_1_port, CARRYB_14_0_port, 
      CARRYB_13_14_port, CARRYB_13_13_port, CARRYB_13_12_port, 
      CARRYB_13_11_port, CARRYB_13_10_port, CARRYB_13_9_port, CARRYB_13_8_port,
      CARRYB_13_7_port, CARRYB_13_6_port, CARRYB_13_5_port, CARRYB_13_4_port, 
      CARRYB_13_3_port, CARRYB_13_2_port, CARRYB_13_1_port, CARRYB_13_0_port, 
      CARRYB_12_14_port, CARRYB_12_13_port, CARRYB_12_12_port, 
      CARRYB_12_11_port, CARRYB_12_10_port, CARRYB_12_9_port, CARRYB_12_8_port,
      CARRYB_12_7_port, CARRYB_12_6_port, CARRYB_12_5_port, CARRYB_12_4_port, 
      CARRYB_12_3_port, CARRYB_12_2_port, CARRYB_12_1_port, CARRYB_12_0_port, 
      CARRYB_11_14_port, CARRYB_11_13_port, CARRYB_11_12_port, 
      CARRYB_11_11_port, CARRYB_11_10_port, CARRYB_11_9_port, CARRYB_11_8_port,
      CARRYB_11_7_port, CARRYB_11_6_port, CARRYB_11_5_port, CARRYB_11_4_port, 
      CARRYB_11_3_port, CARRYB_11_2_port, CARRYB_11_1_port, CARRYB_11_0_port, 
      CARRYB_10_14_port, CARRYB_10_13_port, CARRYB_10_12_port, 
      CARRYB_10_11_port, CARRYB_10_10_port, CARRYB_10_9_port, CARRYB_10_8_port,
      CARRYB_10_7_port, CARRYB_10_6_port, CARRYB_10_5_port, CARRYB_10_4_port, 
      CARRYB_10_3_port, CARRYB_10_2_port, CARRYB_10_1_port, CARRYB_10_0_port, 
      CARRYB_9_14_port, CARRYB_9_13_port, CARRYB_9_12_port, CARRYB_9_11_port, 
      CARRYB_9_10_port, CARRYB_9_9_port, CARRYB_9_8_port, CARRYB_9_7_port, 
      CARRYB_9_6_port, CARRYB_9_5_port, CARRYB_9_4_port, CARRYB_9_3_port, 
      CARRYB_9_2_port, CARRYB_9_1_port, CARRYB_9_0_port, CARRYB_8_14_port, 
      CARRYB_8_13_port, CARRYB_8_12_port, CARRYB_8_11_port, CARRYB_8_10_port, 
      CARRYB_8_9_port, CARRYB_8_8_port, CARRYB_8_7_port, CARRYB_8_6_port, 
      CARRYB_8_5_port, CARRYB_8_4_port, CARRYB_8_3_port, CARRYB_8_2_port, 
      CARRYB_8_1_port, CARRYB_8_0_port, CARRYB_7_14_port, CARRYB_7_13_port, 
      CARRYB_7_12_port, CARRYB_7_11_port, CARRYB_7_10_port, CARRYB_7_9_port, 
      CARRYB_7_8_port, CARRYB_7_7_port, CARRYB_7_6_port, CARRYB_7_5_port, 
      CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, CARRYB_7_1_port, 
      CARRYB_7_0_port, CARRYB_6_14_port, CARRYB_6_13_port, CARRYB_6_12_port, 
      CARRYB_6_11_port, CARRYB_6_10_port, CARRYB_6_9_port, CARRYB_6_8_port, 
      CARRYB_6_7_port, CARRYB_6_6_port, CARRYB_6_5_port, CARRYB_6_3_port, 
      CARRYB_6_2_port, CARRYB_6_1_port, CARRYB_6_0_port, CARRYB_5_14_port, 
      CARRYB_5_13_port, CARRYB_5_12_port, CARRYB_5_11_port, CARRYB_5_10_port, 
      CARRYB_5_9_port, CARRYB_5_8_port, CARRYB_5_7_port, CARRYB_5_6_port, 
      CARRYB_5_5_port, CARRYB_5_4_port, CARRYB_5_3_port, CARRYB_5_2_port, 
      CARRYB_5_1_port, CARRYB_5_0_port, CARRYB_4_14_port, CARRYB_4_13_port, 
      CARRYB_4_12_port, CARRYB_4_11_port, CARRYB_4_10_port, CARRYB_4_9_port, 
      CARRYB_4_8_port, CARRYB_4_7_port, CARRYB_4_6_port, CARRYB_4_5_port, 
      CARRYB_4_3_port, CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, 
      CARRYB_3_14_port, CARRYB_3_13_port, CARRYB_3_12_port, CARRYB_3_11_port, 
      CARRYB_3_10_port, CARRYB_3_9_port, CARRYB_3_8_port, CARRYB_3_7_port, 
      CARRYB_3_6_port, CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, 
      CARRYB_3_2_port, CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_14_port, 
      CARRYB_2_13_port, CARRYB_2_12_port, CARRYB_2_11_port, CARRYB_2_10_port, 
      CARRYB_2_9_port, CARRYB_2_8_port, CARRYB_2_7_port, CARRYB_2_6_port, 
      CARRYB_2_5_port, CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, 
      CARRYB_2_1_port, CARRYB_2_0_port, CARRYB_1_13_port, CARRYB_1_12_port, 
      CARRYB_1_9_port, SUMB_15_15_port, SUMB_15_14_port, SUMB_15_13_port, 
      SUMB_15_12_port, SUMB_15_11_port, SUMB_15_10_port, SUMB_15_9_port, 
      SUMB_15_8_port, SUMB_15_7_port, SUMB_15_6_port, SUMB_15_5_port, 
      SUMB_15_4_port, SUMB_15_3_port, SUMB_15_2_port, SUMB_15_1_port, 
      SUMB_15_0_port, SUMB_14_14_port, SUMB_14_13_port, SUMB_14_12_port, 
      SUMB_14_11_port, SUMB_14_10_port, SUMB_14_9_port, SUMB_14_8_port, 
      SUMB_14_7_port, SUMB_14_6_port, SUMB_14_5_port, SUMB_14_4_port, 
      SUMB_14_3_port, SUMB_14_2_port, SUMB_14_1_port, SUMB_13_14_port, 
      SUMB_13_13_port, SUMB_13_12_port, SUMB_13_11_port, SUMB_13_10_port, 
      SUMB_13_9_port, SUMB_13_8_port, SUMB_13_7_port, SUMB_13_6_port, 
      SUMB_13_5_port, SUMB_13_4_port, SUMB_13_3_port, SUMB_13_2_port, 
      SUMB_13_1_port, SUMB_12_14_port, SUMB_12_13_port, SUMB_12_12_port, 
      SUMB_12_11_port, SUMB_12_10_port, SUMB_12_9_port, SUMB_12_8_port, 
      SUMB_12_7_port, SUMB_12_6_port, SUMB_12_5_port, SUMB_12_4_port, 
      SUMB_12_3_port, SUMB_12_2_port, SUMB_12_1_port, SUMB_11_14_port, 
      SUMB_11_13_port, SUMB_11_12_port, SUMB_11_11_port, SUMB_11_10_port, 
      SUMB_11_9_port, SUMB_11_8_port, SUMB_11_6_port, SUMB_11_5_port, 
      SUMB_11_2_port, SUMB_11_1_port, SUMB_10_14_port, SUMB_10_13_port, 
      SUMB_10_12_port, SUMB_10_11_port, SUMB_10_10_port, SUMB_10_9_port, 
      SUMB_10_8_port, SUMB_10_7_port, SUMB_10_6_port, SUMB_10_5_port, 
      SUMB_10_4_port, SUMB_10_3_port, SUMB_10_2_port, SUMB_10_1_port, 
      SUMB_9_14_port, SUMB_9_13_port, SUMB_9_12_port, SUMB_9_11_port, 
      SUMB_9_10_port, SUMB_9_9_port, SUMB_9_8_port, SUMB_9_7_port, 
      SUMB_9_6_port, SUMB_9_5_port, SUMB_9_4_port, SUMB_9_3_port, SUMB_9_2_port
      , SUMB_9_1_port, SUMB_8_14_port, SUMB_8_13_port, SUMB_8_12_port, 
      SUMB_8_11_port, SUMB_8_10_port, SUMB_8_9_port, SUMB_8_8_port, 
      SUMB_8_7_port, SUMB_8_6_port, SUMB_8_5_port, SUMB_8_4_port, SUMB_8_3_port
      , SUMB_8_2_port, SUMB_8_1_port, SUMB_7_14_port, SUMB_7_13_port, 
      SUMB_7_12_port, SUMB_7_11_port, SUMB_7_10_port, SUMB_7_9_port, 
      SUMB_7_8_port, SUMB_7_7_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port
      , SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_6_14_port, 
      SUMB_6_13_port, SUMB_6_12_port, SUMB_6_11_port, SUMB_6_10_port, 
      SUMB_6_9_port, SUMB_6_8_port, SUMB_6_7_port, SUMB_6_6_port, SUMB_6_5_port
      , SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, SUMB_6_1_port, 
      SUMB_5_14_port, SUMB_5_13_port, SUMB_5_12_port, SUMB_5_11_port, 
      SUMB_5_10_port, SUMB_5_9_port, SUMB_5_8_port, SUMB_5_7_port, 
      SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port, SUMB_5_2_port
      , SUMB_5_1_port, SUMB_4_14_port, SUMB_4_13_port, SUMB_4_12_port, 
      SUMB_4_11_port, SUMB_4_10_port, SUMB_4_9_port, SUMB_4_7_port, 
      SUMB_4_6_port, SUMB_4_5_port, SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port
      , SUMB_4_1_port, SUMB_3_14_port, SUMB_3_13_port, SUMB_3_12_port, 
      SUMB_3_11_port, SUMB_3_10_port, SUMB_3_9_port, SUMB_3_8_port, 
      SUMB_3_7_port, SUMB_3_6_port, SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port
      , SUMB_3_2_port, SUMB_3_1_port, SUMB_2_14_port, SUMB_2_13_port, 
      SUMB_2_12_port, SUMB_2_10_port, SUMB_2_9_port, SUMB_2_8_port, 
      SUMB_2_7_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, SUMB_1_14_port, SUMB_1_13_port, 
      SUMB_1_12_port, SUMB_1_11_port, SUMB_1_10_port, SUMB_1_9_port, 
      SUMB_1_8_port, SUMB_1_7_port, SUMB_1_6_port, SUMB_1_5_port, SUMB_1_4_port
      , SUMB_1_3_port, SUMB_1_2_port, SUMB_1_1_port, A1_28_port, A1_27_port, 
      A1_26_port, A1_25_port, A1_24_port, A1_23_port, A1_22_port, A1_21_port, 
      A1_20_port, A1_19_port, A1_18_port, A1_17_port, A1_16_port, A1_15_port, 
      A1_14_port, A1_13_port, A1_12_port, A1_11_port, A1_10_port, A1_9_port, 
      A1_8_port, A1_7_port, A1_6_port, A1_5_port, A1_4_port, A1_3_port, 
      A1_2_port, A1_1_port, A1_0_port, A2_14_port, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
      n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
      n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
      n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
      n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
      n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
      n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
      n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
      n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
      n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
      n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
      n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
      n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, 
      n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
      n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
      n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
      n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
      n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, 
      n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
      n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, 
      n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, 
      n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, 
      n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, 
      n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, 
      n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, 
      n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
      n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, 
      n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, 
      n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, 
      n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, 
      n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, 
      n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, 
      n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, 
      n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, 
      n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, 
      n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, 
      n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, 
      n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, 
      n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, 
      n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, 
      n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008
      , n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, 
      n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, 
      n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
      n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
      n1049, n1050, n1051, n1052, n1053, n_1195, n_1196, n_1197, n_1198, n_1199
      , n_1200, n_1201, n_1202, n_1203 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_5 : FAX1 port map( A => ab_15_5_port, B => CARRYB_14_5_port, C => 
                           SUMB_14_6_port, YC => CARRYB_15_5_port, YS => 
                           SUMB_15_5_port);
   S4_8 : FAX1 port map( A => ab_15_8_port, B => CARRYB_14_8_port, C => 
                           SUMB_14_9_port, YC => CARRYB_15_8_port, YS => 
                           SUMB_15_8_port);
   S4_9 : FAX1 port map( A => ab_15_9_port, B => CARRYB_14_9_port, C => 
                           SUMB_14_10_port, YC => CARRYB_15_9_port, YS => 
                           SUMB_15_9_port);
   S4_10 : FAX1 port map( A => ab_15_10_port, B => CARRYB_14_10_port, C => 
                           SUMB_14_11_port, YC => CARRYB_15_10_port, YS => 
                           SUMB_15_10_port);
   S4_11 : FAX1 port map( A => ab_15_11_port, B => CARRYB_14_11_port, C => 
                           SUMB_14_12_port, YC => CARRYB_15_11_port, YS => 
                           SUMB_15_11_port);
   S4_12 : FAX1 port map( A => ab_15_12_port, B => CARRYB_14_12_port, C => 
                           SUMB_14_13_port, YC => CARRYB_15_12_port, YS => 
                           SUMB_15_12_port);
   S4_13 : FAX1 port map( A => ab_15_13_port, B => CARRYB_14_13_port, C => 
                           SUMB_14_14_port, YC => CARRYB_15_13_port, YS => 
                           SUMB_15_13_port);
   S5_14 : FAX1 port map( A => ab_15_14_port, B => CARRYB_14_14_port, C => 
                           ab_14_15_port, YC => CARRYB_15_14_port, YS => 
                           SUMB_15_14_port);
   S14_15 : FAX1 port map( A => n1050, B => n1049, C => ab_15_15_port, YC => 
                           CARRYB_15_15_port, YS => SUMB_15_15_port);
   S2_14_9 : FAX1 port map( A => ab_14_9_port, B => CARRYB_13_9_port, C => 
                           SUMB_13_10_port, YC => CARRYB_14_9_port, YS => 
                           SUMB_14_9_port);
   S2_14_10 : FAX1 port map( A => ab_14_10_port, B => CARRYB_13_10_port, C => 
                           SUMB_13_11_port, YC => CARRYB_14_10_port, YS => 
                           SUMB_14_10_port);
   S2_14_11 : FAX1 port map( A => ab_14_11_port, B => CARRYB_13_11_port, C => 
                           SUMB_13_12_port, YC => CARRYB_14_11_port, YS => 
                           SUMB_14_11_port);
   S2_14_12 : FAX1 port map( A => ab_14_12_port, B => CARRYB_13_12_port, C => 
                           SUMB_13_13_port, YC => CARRYB_14_12_port, YS => 
                           SUMB_14_12_port);
   S2_14_13 : FAX1 port map( A => ab_14_13_port, B => CARRYB_13_13_port, C => 
                           SUMB_13_14_port, YC => CARRYB_14_13_port, YS => 
                           SUMB_14_13_port);
   S3_14_14 : FAX1 port map( A => ab_14_14_port, B => CARRYB_13_14_port, C => 
                           ab_13_15_port, YC => CARRYB_14_14_port, YS => 
                           SUMB_14_14_port);
   S2_13_9 : FAX1 port map( A => ab_13_9_port, B => CARRYB_12_9_port, C => 
                           SUMB_12_10_port, YC => CARRYB_13_9_port, YS => 
                           SUMB_13_9_port);
   S2_13_10 : FAX1 port map( A => ab_13_10_port, B => CARRYB_12_10_port, C => 
                           SUMB_12_11_port, YC => CARRYB_13_10_port, YS => 
                           SUMB_13_10_port);
   S2_13_11 : FAX1 port map( A => ab_13_11_port, B => CARRYB_12_11_port, C => 
                           SUMB_12_12_port, YC => CARRYB_13_11_port, YS => 
                           SUMB_13_11_port);
   S2_13_12 : FAX1 port map( A => ab_13_12_port, B => CARRYB_12_12_port, C => 
                           SUMB_12_13_port, YC => CARRYB_13_12_port, YS => 
                           SUMB_13_12_port);
   S2_13_13 : FAX1 port map( A => ab_13_13_port, B => CARRYB_12_13_port, C => 
                           SUMB_12_14_port, YC => CARRYB_13_13_port, YS => 
                           SUMB_13_13_port);
   S3_13_14 : FAX1 port map( A => ab_13_14_port, B => CARRYB_12_14_port, C => 
                           ab_12_15_port, YC => CARRYB_13_14_port, YS => 
                           SUMB_13_14_port);
   S2_12_11 : FAX1 port map( A => ab_12_11_port, B => CARRYB_11_11_port, C => 
                           SUMB_11_12_port, YC => CARRYB_12_11_port, YS => 
                           SUMB_12_11_port);
   S2_12_12 : FAX1 port map( A => ab_12_12_port, B => CARRYB_11_12_port, C => 
                           SUMB_11_13_port, YC => CARRYB_12_12_port, YS => 
                           SUMB_12_12_port);
   S2_12_13 : FAX1 port map( A => ab_12_13_port, B => CARRYB_11_13_port, C => 
                           SUMB_11_14_port, YC => CARRYB_12_13_port, YS => 
                           SUMB_12_13_port);
   S3_12_14 : FAX1 port map( A => ab_12_14_port, B => CARRYB_11_14_port, C => 
                           ab_11_15_port, YC => CARRYB_12_14_port, YS => 
                           SUMB_12_14_port);
   S2_11_9 : FAX1 port map( A => ab_11_9_port, B => CARRYB_10_9_port, C => 
                           SUMB_10_10_port, YC => CARRYB_11_9_port, YS => 
                           SUMB_11_9_port);
   S2_11_11 : FAX1 port map( A => ab_11_11_port, B => CARRYB_10_11_port, C => 
                           SUMB_10_12_port, YC => CARRYB_11_11_port, YS => 
                           SUMB_11_11_port);
   S2_11_12 : FAX1 port map( A => ab_11_12_port, B => CARRYB_10_12_port, C => 
                           SUMB_10_13_port, YC => CARRYB_11_12_port, YS => 
                           SUMB_11_12_port);
   S2_11_13 : FAX1 port map( A => ab_11_13_port, B => CARRYB_10_13_port, C => 
                           SUMB_10_14_port, YC => CARRYB_11_13_port, YS => 
                           SUMB_11_13_port);
   S3_11_14 : FAX1 port map( A => ab_11_14_port, B => CARRYB_10_14_port, C => 
                           ab_10_15_port, YC => CARRYB_11_14_port, YS => 
                           SUMB_11_14_port);
   S2_10_10 : FAX1 port map( A => ab_10_10_port, B => CARRYB_9_10_port, C => 
                           SUMB_9_11_port, YC => CARRYB_10_10_port, YS => 
                           SUMB_10_10_port);
   S2_10_11 : FAX1 port map( A => ab_10_11_port, B => CARRYB_9_11_port, C => 
                           SUMB_9_12_port, YC => CARRYB_10_11_port, YS => 
                           SUMB_10_11_port);
   S2_10_12 : FAX1 port map( A => ab_10_12_port, B => CARRYB_9_12_port, C => 
                           SUMB_9_13_port, YC => CARRYB_10_12_port, YS => 
                           SUMB_10_12_port);
   S2_10_13 : FAX1 port map( A => ab_10_13_port, B => CARRYB_9_13_port, C => 
                           SUMB_9_14_port, YC => CARRYB_10_13_port, YS => 
                           SUMB_10_13_port);
   S3_10_14 : FAX1 port map( A => ab_10_14_port, B => CARRYB_9_14_port, C => 
                           ab_9_15_port, YC => CARRYB_10_14_port, YS => 
                           SUMB_10_14_port);
   S2_9_12 : FAX1 port map( A => ab_9_12_port, B => CARRYB_8_12_port, C => 
                           SUMB_8_13_port, YC => CARRYB_9_12_port, YS => 
                           SUMB_9_12_port);
   S3_9_14 : FAX1 port map( A => ab_9_14_port, B => CARRYB_8_14_port, C => 
                           ab_8_15_port, YC => CARRYB_9_14_port, YS => 
                           SUMB_9_14_port);
   S1_8_0 : FAX1 port map( A => ab_8_0_port, B => CARRYB_7_0_port, C => 
                           SUMB_7_1_port, YC => CARRYB_8_0_port, YS => 
                           A1_6_port);
   S2_8_9 : FAX1 port map( A => ab_8_9_port, B => CARRYB_7_9_port, C => 
                           SUMB_7_10_port, YC => CARRYB_8_9_port, YS => 
                           SUMB_8_9_port);
   S3_8_14 : FAX1 port map( A => ab_8_14_port, B => CARRYB_7_14_port, C => 
                           ab_7_15_port, YC => CARRYB_8_14_port, YS => 
                           SUMB_8_14_port);
   S2_7_1 : FAX1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, C => 
                           SUMB_6_2_port, YC => CARRYB_7_1_port, YS => 
                           SUMB_7_1_port);
   S2_7_13 : FAX1 port map( A => ab_7_13_port, B => CARRYB_6_13_port, C => 
                           SUMB_6_14_port, YC => CARRYB_7_13_port, YS => 
                           SUMB_7_13_port);
   S3_7_14 : FAX1 port map( A => ab_7_14_port, B => CARRYB_6_14_port, C => 
                           ab_6_15_port, YC => CARRYB_7_14_port, YS => 
                           SUMB_7_14_port);
   S1_6_0 : FAX1 port map( A => ab_6_0_port, B => SUMB_5_1_port, C => 
                           CARRYB_5_0_port, YC => CARRYB_6_0_port, YS => 
                           A1_4_port);
   S3_6_14 : FAX1 port map( A => ab_6_14_port, B => CARRYB_5_14_port, C => 
                           ab_5_15_port, YC => CARRYB_6_14_port, YS => 
                           SUMB_6_14_port);
   S1_5_0 : FAX1 port map( A => ab_5_0_port, B => n908, C => SUMB_4_1_port, YC 
                           => CARRYB_5_0_port, YS => A1_3_port);
   S1_4_0 : FAX1 port map( A => ab_4_0_port, B => n906, C => SUMB_3_1_port, YC 
                           => CARRYB_4_0_port, YS => A1_2_port);
   S3_4_14 : FAX1 port map( A => ab_4_14_port, B => CARRYB_3_14_port, C => 
                           ab_3_15_port, YC => CARRYB_4_14_port, YS => 
                           SUMB_4_14_port);
   S1_3_0 : FAX1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, C => 
                           SUMB_2_1_port, YC => CARRYB_3_0_port, YS => 
                           A1_1_port);
   S1_2_0 : FAX1 port map( A => ab_2_0_port, B => n74, C => SUMB_1_1_port, YC 
                           => CARRYB_2_0_port, YS => A1_0_port);
   S2_2_1 : FAX1 port map( A => ab_2_1_port, B => n969, C => SUMB_1_2_port, YC 
                           => CARRYB_2_1_port, YS => SUMB_2_1_port);
   FS_1 : matrix_math_DW01_add_24 port map( A(29) => n1048, A(28) => A1_28_port
                           , A(27) => A1_27_port, A(26) => A1_26_port, A(25) =>
                           A1_25_port, A(24) => A1_24_port, A(23) => A1_23_port
                           , A(22) => A1_22_port, A(21) => A1_21_port, A(20) =>
                           A1_20_port, A(19) => A1_19_port, A(18) => A1_18_port
                           , A(17) => A1_17_port, A(16) => A1_16_port, A(15) =>
                           A1_15_port, A(14) => A1_14_port, A(13) => A1_13_port
                           , A(12) => A1_12_port, A(11) => A1_11_port, A(10) =>
                           A1_10_port, A(9) => A1_9_port, A(8) => A1_8_port, 
                           A(7) => A1_7_port, A(6) => A1_6_port, A(5) => 
                           A1_5_port, A(4) => A1_4_port, A(3) => A1_3_port, 
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(29) => n73, B(28) => n72, B(27) => n71,
                           B(26) => n70, B(25) => n69, B(24) => n68, B(23) => 
                           n67, B(22) => n66, B(21) => n80, B(20) => n973, 
                           B(19) => n968, B(18) => n967, B(17) => n966, B(16) 
                           => n971, B(15) => n972, B(14) => A2_14_port, B(13) 
                           => n1053, B(12) => n1053, B(11) => n1053, B(10) => 
                           n1053, B(9) => n1053, B(8) => n1053, B(7) => n1053, 
                           B(6) => n1053, B(5) => n1053, B(4) => n1053, B(3) =>
                           n1053, B(2) => n1053, B(1) => n1053, B(0) => 
                           X_Logic0_port, CI => X_Logic0_port, SUM(29) => 
                           n_1195, SUM(28) => n_1196, SUM(27) => n_1197, 
                           SUM(26) => n_1198, SUM(25) => n_1199, SUM(24) => 
                           n_1200, SUM(23) => n_1201, SUM(22) => n_1202, 
                           SUM(21) => PRODUCT(23), SUM(20) => PRODUCT(22), 
                           SUM(19) => PRODUCT(21), SUM(18) => PRODUCT(20), 
                           SUM(17) => PRODUCT(19), SUM(16) => PRODUCT(18), 
                           SUM(15) => PRODUCT(17), SUM(14) => PRODUCT(16), 
                           SUM(13) => PRODUCT(15), SUM(12) => PRODUCT(14), 
                           SUM(11) => PRODUCT(13), SUM(10) => PRODUCT(12), 
                           SUM(9) => PRODUCT(11), SUM(8) => PRODUCT(10), SUM(7)
                           => PRODUCT(9), SUM(6) => PRODUCT(8), SUM(5) => 
                           PRODUCT(7), SUM(4) => PRODUCT(6), SUM(3) => 
                           PRODUCT(5), SUM(2) => PRODUCT(4), SUM(1) => 
                           PRODUCT(3), SUM(0) => PRODUCT(2), CO => n_1203);
   U2 : XOR2X1 port map( A => n14, B => n3, Y => SUMB_9_5_port);
   U3 : XNOR2X1 port map( A => n129, B => n130, Y => n3);
   U4 : XOR2X1 port map( A => n4, B => n146, Y => SUMB_10_5_port);
   U5 : XNOR2X1 port map( A => CARRYB_9_5_port, B => n157, Y => n4);
   U6 : BUFX2 port map( A => n76, Y => n5);
   U7 : XNOR2X1 port map( A => n6, B => SUMB_4_10_port, Y => SUMB_5_9_port);
   U8 : XNOR2X1 port map( A => CARRYB_4_9_port, B => ab_5_9_port, Y => n6);
   U9 : XNOR2X1 port map( A => n7, B => SUMB_5_9_port, Y => SUMB_6_8_port);
   U10 : XOR2X1 port map( A => CARRYB_5_8_port, B => n175, Y => n7);
   U11 : XNOR2X1 port map( A => n8, B => n297, Y => n223);
   U12 : XOR2X1 port map( A => n222, B => n82, Y => n8);
   U13 : INVX2 port map( A => n763, Y => n9);
   U14 : INVX2 port map( A => n9, Y => n10);
   U15 : BUFX2 port map( A => n606, Y => n11);
   U16 : BUFX2 port map( A => n639, Y => n12);
   U17 : INVX2 port map( A => SUMB_9_9_port, Y => n59);
   U18 : BUFX2 port map( A => n765, Y => n13);
   U19 : XOR2X1 port map( A => CARRYB_8_5_port, B => n224, Y => n14);
   U20 : BUFX2 port map( A => CARRYB_5_3_port, Y => n15);
   U21 : NAND3X1 port map( A => n735, B => n734, C => n733, Y => n16);
   U22 : INVX2 port map( A => SUMB_12_2_port, Y => n320);
   U23 : XNOR2X1 port map( A => n17, B => SUMB_14_1_port, Y => SUMB_15_0_port);
   U24 : XNOR2X1 port map( A => CARRYB_14_0_port, B => n50, Y => n17);
   U25 : XNOR2X1 port map( A => n18, B => n253, Y => SUMB_9_4_port);
   U26 : XOR2X1 port map( A => CARRYB_8_4_port, B => ab_9_4_port, Y => n18);
   U27 : BUFX2 port map( A => CARRYB_12_7_port, Y => n19);
   U28 : XOR2X1 port map( A => SUMB_8_7_port, B => n20, Y => SUMB_9_6_port);
   U29 : XOR2X1 port map( A => CARRYB_8_6_port, B => ab_9_6_port, Y => n20);
   U30 : BUFX2 port map( A => SUMB_15_3_port, Y => n21);
   U31 : AND2X2 port map( A => CARRYB_15_2_port, B => n21, Y => n966);
   U32 : XOR2X1 port map( A => n22, B => SUMB_8_8_port, Y => SUMB_9_7_port);
   U33 : XOR2X1 port map( A => CARRYB_8_7_port, B => ab_9_7_port, Y => n22);
   U34 : XOR2X1 port map( A => n23, B => n5, Y => SUMB_12_6_port);
   U35 : XNOR2X1 port map( A => CARRYB_11_6_port, B => n244, Y => n23);
   U36 : BUFX2 port map( A => n898, Y => n24);
   U37 : XOR2X1 port map( A => CARRYB_11_4_port, B => n25, Y => n339);
   U38 : INVX8 port map( A => ab_12_4_port, Y => n25);
   U39 : BUFX2 port map( A => CARRYB_7_11_port, Y => n26);
   U40 : INVX2 port map( A => SUMB_7_7_port, Y => n130);
   U41 : XOR2X1 port map( A => n86, B => n27, Y => SUMB_14_4_port);
   U42 : XNOR2X1 port map( A => CARRYB_13_4_port, B => ab_14_4_port, Y => n27);
   U43 : XNOR2X1 port map( A => n28, B => SUMB_12_6_port, Y => SUMB_13_5_port);
   U44 : XNOR2X1 port map( A => CARRYB_12_5_port, B => ab_13_5_port, Y => n28);
   U45 : XOR2X1 port map( A => n976, B => n29, Y => SUMB_2_13_port);
   U46 : XNOR2X1 port map( A => SUMB_1_14_port, B => ab_2_13_port, Y => n29);
   U47 : XNOR2X1 port map( A => n30, B => SUMB_6_9_port, Y => SUMB_7_8_port);
   U48 : XNOR2X1 port map( A => CARRYB_6_8_port, B => ab_7_8_port, Y => n30);
   U49 : XOR2X1 port map( A => n158, B => n31, Y => n32);
   U50 : NAND2X1 port map( A => n206, B => n1007, Y => n31);
   U51 : XNOR2X1 port map( A => n32, B => n271, Y => SUMB_2_8_port);
   U52 : BUFX2 port map( A => n883, Y => n33);
   U53 : XNOR2X1 port map( A => CARRYB_14_4_port, B => n34, Y => n676);
   U54 : INVX8 port map( A => ab_15_4_port, Y => n34);
   U55 : INVX1 port map( A => SUMB_13_1_port, Y => n35);
   U56 : INVX1 port map( A => n35, Y => n36);
   U57 : XOR2X1 port map( A => CARRYB_7_4_port, B => n321, Y => n410);
   U58 : XOR2X1 port map( A => n489, B => n37, Y => n267);
   U59 : INVX8 port map( A => n65, Y => n37);
   U60 : NAND3X1 port map( A => n837, B => n839, C => n838, Y => n38);
   U61 : XOR2X1 port map( A => n39, B => n542, Y => SUMB_7_6_port);
   U62 : XNOR2X1 port map( A => CARRYB_6_6_port, B => ab_7_6_port, Y => n39);
   U63 : INVX1 port map( A => n1023, Y => n40);
   U64 : INVX2 port map( A => n1022, Y => n1023);
   U65 : AND2X2 port map( A => n810, B => n812, Y => n79);
   U66 : AND2X1 port map( A => n236, B => n993, Y => ab_2_1_port);
   U67 : AND2X2 port map( A => n206, B => n1007, Y => n41);
   U68 : XOR2X1 port map( A => SUMB_11_1_port, B => ab_12_0_port, Y => n42);
   U69 : XOR2X1 port map( A => CARRYB_11_0_port, B => n42, Y => A1_10_port);
   U70 : NAND2X1 port map( A => CARRYB_11_0_port, B => SUMB_11_1_port, Y => n43
                           );
   U71 : NAND2X1 port map( A => CARRYB_11_0_port, B => ab_12_0_port, Y => n44);
   U72 : NAND2X1 port map( A => SUMB_11_1_port, B => ab_12_0_port, Y => n45);
   U73 : NAND3X1 port map( A => n44, B => n43, C => n45, Y => CARRYB_12_0_port)
                           ;
   U74 : XOR2X1 port map( A => CARRYB_3_7_port, B => n46, Y => n532);
   U75 : INVX8 port map( A => ab_4_7_port, Y => n46);
   U76 : XOR2X1 port map( A => n47, B => n233, Y => SUMB_6_4_port);
   U77 : INVX2 port map( A => n47, Y => n48);
   U78 : INVX2 port map( A => n431, Y => n47);
   U79 : INVX2 port map( A => SUMB_8_5_port, Y => n253);
   U80 : XNOR2X1 port map( A => n49, B => SUMB_9_7_port, Y => SUMB_10_6_port);
   U81 : XNOR2X1 port map( A => CARRYB_9_6_port, B => ab_10_6_port, Y => n49);
   U82 : INVX8 port map( A => n52, Y => n50);
   U83 : INVX2 port map( A => n1010, Y => n51);
   U84 : INVX2 port map( A => B(10), Y => n1010);
   U85 : INVX8 port map( A => ab_15_0_port, Y => n52);
   U86 : NAND3X1 port map( A => n767, B => n768, C => n769, Y => n53);
   U87 : XOR2X1 port map( A => n54, B => n55, Y => SUMB_4_6_port);
   U88 : XNOR2X1 port map( A => CARRYB_3_6_port, B => ab_4_6_port, Y => n54);
   U89 : INVX1 port map( A => SUMB_3_7_port, Y => n55);
   U90 : NAND3X1 port map( A => n730, B => n731, C => n732, Y => n56);
   U91 : BUFX2 port map( A => SUMB_7_9_port, Y => n57);
   U92 : XOR2X1 port map( A => n58, B => n59, Y => SUMB_10_8_port);
   U93 : XNOR2X1 port map( A => CARRYB_9_8_port, B => ab_10_8_port, Y => n58);
   U94 : NAND3X1 port map( A => n309, B => n308, C => n310, Y => n60);
   U95 : INVX4 port map( A => n996, Y => n983);
   U96 : INVX4 port map( A => B(3), Y => n996);
   U97 : INVX1 port map( A => B(6), Y => n1002);
   U98 : AND2X2 port map( A => n439, B => ab_0_8_port, Y => n61);
   U99 : INVX4 port map( A => n1004, Y => n1005);
   U100 : INVX4 port map( A => n1010, Y => n1011);
   U101 : NOR2X1 port map( A => n1000, B => n40, Y => n62);
   U102 : AND2X2 port map( A => ab_0_3_port, B => n964, Y => n63);
   U103 : XNOR2X1 port map( A => CARRYB_14_1_port, B => n64, Y => n561);
   U104 : INVX8 port map( A => ab_15_1_port, Y => n64);
   U105 : INVX1 port map( A => CARRYB_8_6_port, Y => n441);
   U106 : INVX8 port map( A => ab_14_3_port, Y => n65);
   U107 : INVX2 port map( A => ab_10_5_port, Y => n157);
   U108 : INVX2 port map( A => ab_11_4_port, Y => n301);
   U109 : INVX2 port map( A => ab_4_9_port, Y => n401);
   U110 : INVX2 port map( A => ab_12_3_port, Y => n149);
   U111 : INVX2 port map( A => ab_6_7_port, Y => n205);
   U112 : INVX2 port map( A => ab_5_7_port, Y => n261);
   U113 : INVX2 port map( A => ab_7_7_port, Y => n440);
   U114 : INVX2 port map( A => ab_12_6_port, Y => n244);
   U115 : INVX2 port map( A => ab_7_10_port, Y => n248);
   U116 : INVX2 port map( A => ab_11_5_port, Y => n298);
   U117 : INVX2 port map( A => ab_10_4_port, Y => n163);
   U118 : INVX2 port map( A => ab_13_2_port, Y => n251);
   U119 : INVX2 port map( A => ab_14_6_port, Y => n186);
   U120 : INVX2 port map( A => ab_6_9_port, Y => n138);
   U121 : INVX2 port map( A => ab_6_8_port, Y => n175);
   U122 : INVX2 port map( A => ab_4_5_port, Y => n182);
   U123 : INVX2 port map( A => ab_7_5_port, Y => n503);
   U124 : INVX2 port map( A => ab_9_5_port, Y => n224);
   U125 : INVX2 port map( A => ab_8_3_port, Y => n755);
   U126 : INVX2 port map( A => ab_8_4_port, Y => n321);
   U127 : INVX2 port map( A => ab_9_9_port, Y => n189);
   U128 : INVX4 port map( A => n1002, Y => n1003);
   U129 : INVX2 port map( A => ab_14_1_port, Y => n530);
   U130 : INVX2 port map( A => n318, Y => n317);
   U131 : INVX2 port map( A => ab_13_8_port, Y => n324);
   U132 : AND2X1 port map( A => SUMB_15_8_port, B => CARRYB_15_7_port, Y => n66
                           );
   U133 : AND2X2 port map( A => SUMB_15_9_port, B => CARRYB_15_8_port, Y => n67
                           );
   U134 : AND2X2 port map( A => SUMB_15_10_port, B => CARRYB_15_9_port, Y => 
                           n68);
   U135 : AND2X2 port map( A => SUMB_15_11_port, B => CARRYB_15_10_port, Y => 
                           n69);
   U136 : AND2X2 port map( A => SUMB_15_12_port, B => CARRYB_15_11_port, Y => 
                           n70);
   U137 : AND2X2 port map( A => SUMB_15_13_port, B => CARRYB_15_12_port, Y => 
                           n71);
   U138 : AND2X2 port map( A => SUMB_15_14_port, B => CARRYB_15_13_port, Y => 
                           n72);
   U139 : AND2X2 port map( A => SUMB_15_15_port, B => CARRYB_15_14_port, Y => 
                           n73);
   U140 : AND2X2 port map( A => ab_0_1_port, B => ab_1_0_port, Y => n74);
   U141 : AND2X2 port map( A => ab_0_15_port, B => ab_1_14_port, Y => n75);
   U142 : XOR2X1 port map( A => SUMB_10_8_port, B => n586, Y => n76);
   U143 : AND2X2 port map( A => ab_0_11_port, B => ab_1_10_port, Y => n77);
   U144 : AND2X2 port map( A => n527, B => n529, Y => n78);
   U145 : AND2X2 port map( A => SUMB_15_7_port, B => CARRYB_15_6_port, Y => n80
                           );
   U146 : XNOR2X1 port map( A => n81, B => SUMB_2_10_port, Y => SUMB_3_9_port);
   U147 : XNOR2X1 port map( A => CARRYB_2_9_port, B => ab_3_9_port, Y => n81);
   U148 : AND2X2 port map( A => n236, B => n1013, Y => n82);
   U149 : XNOR2X1 port map( A => ab_0_10_port, B => n83, Y => SUMB_1_9_port);
   U150 : NAND2X1 port map( A => B(9), B => n322, Y => n83);
   U151 : NAND3X1 port map( A => n887, B => n888, C => n889, Y => n84);
   U152 : NAND3X1 port map( A => n404, B => n403, C => n405, Y => n85);
   U153 : INVX2 port map( A => CARRYB_15_5_port, Y => n318);
   U154 : INVX1 port map( A => SUMB_13_5_port, Y => n86);
   U155 : NAND3X1 port map( A => n714, B => n715, C => n716, Y => n87);
   U156 : BUFX2 port map( A => n638, Y => n88);
   U157 : BUFX2 port map( A => SUMB_9_1_port, Y => n89);
   U158 : XOR2X1 port map( A => n90, B => n272, Y => SUMB_6_7_port);
   U159 : XOR2X1 port map( A => SUMB_5_8_port, B => n205, Y => n90);
   U160 : NAND3X1 port map( A => n679, B => n678, C => n677, Y => 
                           CARRYB_15_4_port);
   U161 : XOR2X1 port map( A => n91, B => n57, Y => SUMB_8_8_port);
   U162 : XOR2X1 port map( A => CARRYB_7_8_port, B => ab_8_8_port, Y => n91);
   U163 : BUFX2 port map( A => CARRYB_7_2_port, Y => n92);
   U164 : XOR2X1 port map( A => n311, B => n312, Y => n93);
   U165 : INVX2 port map( A => SUMB_10_5_port, Y => n311);
   U166 : BUFX2 port map( A => CARRYB_3_10_port, Y => n94);
   U167 : XOR2X1 port map( A => n152, B => n128, Y => n95);
   U168 : BUFX2 port map( A => CARRYB_3_5_port, Y => n96);
   U169 : XOR2X1 port map( A => n172, B => n215, Y => n97);
   U170 : NAND3X1 port map( A => n675, B => n673, C => n674, Y => n98);
   U171 : NAND3X1 port map( A => n778, B => n779, C => n780, Y => n99);
   U172 : XOR2X1 port map( A => n410, B => n534, Y => n100);
   U173 : INVX2 port map( A => SUMB_7_5_port, Y => n534);
   U174 : XOR2X1 port map( A => CARRYB_9_3_port, B => ab_10_3_port, Y => n449);
   U175 : AND2X2 port map( A => ab_1_8_port, B => ab_0_9_port, Y => n737);
   U176 : XOR2X1 port map( A => CARRYB_5_13_port, B => ab_6_13_port, Y => n101)
                           ;
   U177 : XOR2X1 port map( A => SUMB_5_14_port, B => n101, Y => SUMB_6_13_port)
                           ;
   U178 : NAND2X1 port map( A => SUMB_5_14_port, B => CARRYB_5_13_port, Y => 
                           n102);
   U179 : NAND2X1 port map( A => SUMB_5_14_port, B => ab_6_13_port, Y => n103);
   U180 : NAND2X1 port map( A => CARRYB_5_13_port, B => ab_6_13_port, Y => n104
                           );
   U181 : NAND3X1 port map( A => n103, B => n102, C => n104, Y => 
                           CARRYB_6_13_port);
   U182 : XOR2X1 port map( A => ab_5_14_port, B => ab_4_15_port, Y => n105);
   U183 : XOR2X1 port map( A => CARRYB_4_14_port, B => n105, Y => 
                           SUMB_5_14_port);
   U184 : NAND2X1 port map( A => CARRYB_4_14_port, B => ab_5_14_port, Y => n106
                           );
   U185 : NAND2X1 port map( A => CARRYB_4_14_port, B => ab_4_15_port, Y => n107
                           );
   U186 : NAND2X1 port map( A => ab_5_14_port, B => ab_4_15_port, Y => n108);
   U187 : NAND3X1 port map( A => n107, B => n106, C => n108, Y => 
                           CARRYB_5_14_port);
   U188 : XOR2X1 port map( A => CARRYB_13_8_port, B => ab_14_8_port, Y => n109)
                           ;
   U189 : XOR2X1 port map( A => SUMB_13_9_port, B => n109, Y => SUMB_14_8_port)
                           ;
   U190 : NAND2X1 port map( A => SUMB_13_9_port, B => CARRYB_13_8_port, Y => 
                           n110);
   U191 : NAND2X1 port map( A => SUMB_13_9_port, B => ab_14_8_port, Y => n111);
   U192 : NAND2X1 port map( A => CARRYB_13_8_port, B => ab_14_8_port, Y => n112
                           );
   U193 : NAND3X1 port map( A => n111, B => n110, C => n112, Y => 
                           CARRYB_14_8_port);
   U194 : XOR2X1 port map( A => CARRYB_10_10_port, B => ab_11_10_port, Y => 
                           n113);
   U195 : XOR2X1 port map( A => SUMB_10_11_port, B => n113, Y => 
                           SUMB_11_10_port);
   U196 : NAND2X1 port map( A => SUMB_10_11_port, B => CARRYB_10_10_port, Y => 
                           n114);
   U197 : NAND2X1 port map( A => SUMB_10_11_port, B => ab_11_10_port, Y => n115
                           );
   U198 : NAND2X1 port map( A => CARRYB_10_10_port, B => ab_11_10_port, Y => 
                           n116);
   U199 : NAND3X1 port map( A => n115, B => n114, C => n116, Y => 
                           CARRYB_11_10_port);
   U200 : BUFX2 port map( A => SUMB_6_12_port, Y => n117);
   U201 : XNOR2X1 port map( A => n118, B => SUMB_5_13_port, Y => SUMB_6_12_port
                           );
   U202 : XOR2X1 port map( A => n711, B => ab_6_12_port, Y => n118);
   U203 : XOR2X1 port map( A => SUMB_15_5_port, B => CARRYB_15_4_port, Y => 
                           A1_18_port);
   U204 : BUFX2 port map( A => n748, Y => n119);
   U205 : BUFX2 port map( A => n794, Y => n120);
   U206 : BUFX2 port map( A => SUMB_4_5_port, Y => n121);
   U207 : NAND3X1 port map( A => n666, B => n664, C => n665, Y => n122);
   U208 : XOR2X1 port map( A => CARRYB_10_7_port, B => ab_11_7_port, Y => n586)
                           ;
   U209 : XOR2X1 port map( A => CARRYB_12_6_port, B => ab_13_6_port, Y => n424)
                           ;
   U210 : BUFX2 port map( A => n698, Y => n123);
   U211 : NAND3X1 port map( A => n587, B => n588, C => n589, Y => n124);
   U212 : XNOR2X1 port map( A => n125, B => SUMB_12_8_port, Y => SUMB_13_7_port
                           );
   U213 : XNOR2X1 port map( A => ab_13_7_port, B => CARRYB_12_7_port, Y => n125
                           );
   U214 : NAND3X1 port map( A => n667, B => n668, C => n669, Y => n126);
   U215 : XOR2X1 port map( A => SUMB_8_9_port, B => n127, Y => SUMB_9_8_port);
   U216 : XOR2X1 port map( A => CARRYB_8_8_port, B => ab_9_8_port, Y => n127);
   U217 : XOR2X1 port map( A => n152, B => n128, Y => SUMB_5_11_port);
   U218 : XOR2X1 port map( A => CARRYB_4_11_port, B => ab_5_11_port, Y => n128)
                           ;
   U219 : XOR2X1 port map( A => n129, B => n130, Y => SUMB_8_6_port);
   U220 : XNOR2X1 port map( A => n147, B => ab_8_6_port, Y => n129);
   U221 : INVX1 port map( A => n1007, Y => n131);
   U222 : INVX4 port map( A => n131, Y => n132);
   U223 : INVX4 port map( A => n1006, Y => n1007);
   U224 : INVX2 port map( A => B(8), Y => n1006);
   U225 : XOR2X1 port map( A => SUMB_11_2_port, B => ab_12_1_port, Y => n169);
   U226 : XNOR2X1 port map( A => n133, B => n100, Y => SUMB_9_3_port);
   U227 : XNOR2X1 port map( A => CARRYB_8_3_port, B => ab_9_3_port, Y => n133);
   U228 : XNOR2X1 port map( A => n134, B => n135, Y => SUMB_11_2_port);
   U229 : XOR2X1 port map( A => CARRYB_10_2_port, B => ab_11_2_port, Y => n134)
                           ;
   U230 : XOR2X1 port map( A => n449, B => n377, Y => n135);
   U231 : INVX2 port map( A => SUMB_6_7_port, Y => n542);
   U232 : XNOR2X1 port map( A => n136, B => SUMB_12_3_port, Y => SUMB_13_2_port
                           );
   U233 : XOR2X1 port map( A => CARRYB_12_2_port, B => n251, Y => n136);
   U234 : XNOR2X1 port map( A => ab_1_11_port, B => n137, Y => SUMB_1_11_port);
   U235 : NAND2X1 port map( A => n266, B => n1015, Y => n137);
   U236 : XNOR2X1 port map( A => n336, B => n138, Y => n726);
   U237 : INVX1 port map( A => SUMB_5_5_port, Y => n431);
   U238 : INVX1 port map( A => n974, Y => CARRYB_1_9_port);
   U239 : XNOR2X1 port map( A => n725, B => n139, Y => SUMB_5_10_port);
   U240 : INVX2 port map( A => SUMB_4_11_port, Y => n139);
   U241 : AND2X1 port map( A => SUMB_15_4_port, B => CARRYB_15_3_port, Y => 
                           n967);
   U242 : XOR2X1 port map( A => SUMB_1_5_port, B => ab_2_4_port, Y => n140);
   U243 : XOR2X1 port map( A => n965, B => n140, Y => SUMB_2_4_port);
   U244 : NAND2X1 port map( A => n965, B => SUMB_1_5_port, Y => n141);
   U245 : NAND2X1 port map( A => n965, B => ab_2_4_port, Y => n142);
   U246 : NAND2X1 port map( A => SUMB_1_5_port, B => ab_2_4_port, Y => n143);
   U247 : NAND3X1 port map( A => n142, B => n141, C => n143, Y => 
                           CARRYB_2_4_port);
   U248 : BUFX2 port map( A => CARRYB_12_0_port, Y => n144);
   U249 : NAND3X1 port map( A => n870, B => n869, C => n871, Y => n145);
   U250 : BUFX2 port map( A => SUMB_9_6_port, Y => n146);
   U251 : NAND3X1 port map( A => n944, B => n943, C => n942, Y => n147);
   U252 : INVX1 port map( A => SUMB_5_10_port, Y => n300);
   U253 : AND2X2 port map( A => n266, B => n1015, Y => n148);
   U254 : XOR2X1 port map( A => CARRYB_11_3_port, B => n149, Y => n195);
   U255 : INVX2 port map( A => n1022, Y => n235);
   U256 : INVX2 port map( A => n1022, Y => n236);
   U257 : INVX1 port map( A => SUMB_1_14_port, Y => n150);
   U258 : INVX1 port map( A => n150, Y => n151);
   U259 : BUFX2 port map( A => SUMB_4_12_port, Y => n152);
   U260 : XOR2X1 port map( A => SUMB_8_11_port, B => ab_9_10_port, Y => n153);
   U261 : XOR2X1 port map( A => n153, B => CARRYB_8_10_port, Y => 
                           SUMB_9_10_port);
   U262 : NAND2X1 port map( A => CARRYB_8_10_port, B => SUMB_8_11_port, Y => 
                           n154);
   U263 : NAND2X1 port map( A => CARRYB_8_10_port, B => ab_9_10_port, Y => n155
                           );
   U264 : NAND2X1 port map( A => SUMB_8_11_port, B => ab_9_10_port, Y => n156);
   U265 : NAND3X1 port map( A => n155, B => n154, C => n156, Y => 
                           CARRYB_9_10_port);
   U266 : INVX1 port map( A => n472, Y => n473);
   U267 : INVX2 port map( A => SUMB_1_9_port, Y => n271);
   U268 : NAND2X1 port map( A => ab_1_8_port, B => ab_0_9_port, Y => n158);
   U269 : XOR2X1 port map( A => n159, B => n160, Y => SUMB_6_1_port);
   U270 : XNOR2X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, Y => n159);
   U271 : INVX1 port map( A => SUMB_5_2_port, Y => n160);
   U272 : XNOR2X1 port map( A => n791, B => n161, Y => SUMB_7_9_port);
   U273 : INVX2 port map( A => SUMB_6_10_port, Y => n161);
   U274 : AND2X2 port map( A => CARRYB_15_1_port, B => SUMB_15_2_port, Y => 
                           n971);
   U275 : BUFX2 port map( A => n835, Y => n162);
   U276 : XOR2X1 port map( A => CARRYB_9_4_port, B => n163, Y => n376);
   U277 : BUFX2 port map( A => SUMB_8_1_port, Y => n164);
   U278 : XOR2X1 port map( A => CARRYB_10_1_port, B => ab_11_1_port, Y => n165)
                           ;
   U279 : XOR2X1 port map( A => n165, B => SUMB_10_2_port, Y => SUMB_11_1_port)
                           ;
   U280 : XNOR2X1 port map( A => n166, B => SUMB_14_3_port, Y => SUMB_15_2_port
                           );
   U281 : XNOR2X1 port map( A => CARRYB_14_2_port, B => ab_15_2_port, Y => n166
                           );
   U282 : XOR2X1 port map( A => n167, B => SUMB_13_7_port, Y => SUMB_14_6_port)
                           ;
   U283 : XNOR2X1 port map( A => CARRYB_13_6_port, B => n186, Y => n167);
   U284 : XNOR2X1 port map( A => n168, B => n171, Y => SUMB_7_5_port);
   U285 : XOR2X1 port map( A => SUMB_6_6_port, B => n503, Y => n168);
   U286 : XNOR2X1 port map( A => n169, B => n170, Y => SUMB_12_1_port);
   U287 : INVX1 port map( A => CARRYB_11_1_port, Y => n170);
   U288 : BUFX2 port map( A => CARRYB_6_5_port, Y => n171);
   U289 : XOR2X1 port map( A => n172, B => n215, Y => SUMB_2_7_port);
   U290 : XNOR2X1 port map( A => n435, B => n314, Y => n172);
   U291 : INVX1 port map( A => CARRYB_2_8_port, Y => n436);
   U292 : NAND3X1 port map( A => n803, B => n802, C => n801, Y => n173);
   U293 : NAND3X1 port map( A => n885, B => n884, C => n886, Y => n174);
   U294 : XNOR2X1 port map( A => n176, B => SUMB_7_8_port, Y => SUMB_8_7_port);
   U295 : XNOR2X1 port map( A => CARRYB_7_7_port, B => ab_8_7_port, Y => n176);
   U296 : XNOR2X1 port map( A => n177, B => n223, Y => SUMB_3_10_port);
   U297 : XNOR2X1 port map( A => CARRYB_2_10_port, B => ab_3_10_port, Y => n177
                           );
   U298 : INVX2 port map( A => n998, Y => n984);
   U299 : INVX4 port map( A => n986, Y => n514);
   U300 : XOR2X1 port map( A => n178, B => CARRYB_5_2_port, Y => SUMB_6_2_port)
                           ;
   U301 : XOR2X1 port map( A => SUMB_5_3_port, B => ab_6_2_port, Y => n178);
   U302 : NAND3X1 port map( A => n257, B => n258, C => n259, Y => n179);
   U303 : NAND3X1 port map( A => n383, B => n382, C => n384, Y => n180);
   U304 : AND2X2 port map( A => ab_0_7_port, B => ab_1_6_port, Y => n181);
   U305 : AND2X2 port map( A => B(6), B => n987, Y => n524);
   U306 : XOR2X1 port map( A => SUMB_3_6_port, B => n182, Y => n234);
   U307 : XOR2X1 port map( A => n183, B => n97, Y => SUMB_3_6_port);
   U308 : XNOR2X1 port map( A => n847, B => ab_3_6_port, Y => n183);
   U309 : XOR2X1 port map( A => CARRYB_7_3_port, B => n755, Y => n216);
   U310 : AND2X2 port map( A => B(9), B => n322, Y => n184);
   U311 : BUFX2 port map( A => CARRYB_4_3_port, Y => n185);
   U312 : BUFX2 port map( A => n894, Y => n187);
   U313 : INVX2 port map( A => SUMB_8_3_port, Y => n608);
   U314 : XOR2X1 port map( A => n448, B => n188, Y => SUMB_8_5_port);
   U315 : INVX2 port map( A => SUMB_7_6_port, Y => n188);
   U316 : XOR2X1 port map( A => n189, B => n220, Y => n194);
   U317 : INVX1 port map( A => n220, Y => n221);
   U318 : NAND3X1 port map( A => n955, B => n954, C => n956, Y => n190);
   U319 : XNOR2X1 port map( A => n191, B => n192, Y => SUMB_7_3_port);
   U320 : XOR2X1 port map( A => n413, B => ab_7_3_port, Y => n191);
   U321 : XOR2X1 port map( A => n233, B => n48, Y => n192);
   U322 : NAND3X1 port map( A => n479, B => n478, C => n480, Y => n193);
   U323 : INVX1 port map( A => CARRYB_6_2_port, Y => n960);
   U324 : XOR2X1 port map( A => n194, B => SUMB_8_10_port, Y => SUMB_9_9_port);
   U325 : XNOR2X1 port map( A => n195, B => n93, Y => SUMB_12_3_port);
   U326 : BUFX2 port map( A => SUMB_3_5_port, Y => n196);
   U327 : NAND3X1 port map( A => n958, B => n959, C => n957, Y => n197);
   U328 : XOR2X1 port map( A => SUMB_3_11_port, B => ab_4_10_port, Y => n198);
   U329 : XOR2X1 port map( A => n94, B => n198, Y => SUMB_4_10_port);
   U330 : NAND2X1 port map( A => SUMB_3_11_port, B => CARRYB_3_10_port, Y => 
                           n199);
   U331 : NAND2X1 port map( A => CARRYB_3_10_port, B => ab_4_10_port, Y => n200
                           );
   U332 : NAND2X1 port map( A => SUMB_3_11_port, B => ab_4_10_port, Y => n201);
   U333 : NAND3X1 port map( A => n200, B => n199, C => n201, Y => 
                           CARRYB_4_10_port);
   U334 : NAND3X1 port map( A => n624, B => n625, C => n626, Y => n202);
   U335 : NAND3X1 port map( A => n764, B => n13, C => n766, Y => n203);
   U336 : NAND3X1 port map( A => n834, B => n836, C => n162, Y => n204);
   U337 : INVX2 port map( A => n1022, Y => n206);
   U338 : XOR2X1 port map( A => n207, B => n208, Y => SUMB_7_4_port);
   U339 : XNOR2X1 port map( A => n122, B => ab_7_4_port, Y => n207);
   U340 : INVX2 port map( A => SUMB_6_5_port, Y => n208);
   U341 : XOR2X1 port map( A => SUMB_3_14_port, B => ab_4_13_port, Y => n209);
   U342 : XOR2X1 port map( A => CARRYB_3_13_port, B => n209, Y => 
                           SUMB_4_13_port);
   U343 : NAND2X1 port map( A => CARRYB_3_13_port, B => SUMB_3_14_port, Y => 
                           n210);
   U344 : NAND2X1 port map( A => CARRYB_3_13_port, B => ab_4_13_port, Y => n211
                           );
   U345 : NAND2X1 port map( A => SUMB_3_14_port, B => ab_4_13_port, Y => n212);
   U346 : NAND3X1 port map( A => n211, B => n210, C => n212, Y => 
                           CARRYB_4_13_port);
   U347 : NAND3X1 port map( A => n391, B => n390, C => n392, Y => n213);
   U348 : INVX1 port map( A => n847, Y => n848);
   U349 : INVX1 port map( A => SUMB_1_12_port, Y => n297);
   U350 : XOR2X1 port map( A => n219, B => n269, Y => n214);
   U351 : BUFX2 port map( A => SUMB_1_8_port, Y => n215);
   U352 : XOR2X1 port map( A => n216, B => n375, Y => SUMB_8_3_port);
   U353 : XNOR2X1 port map( A => n519, B => n217, Y => SUMB_2_6_port);
   U354 : INVX1 port map( A => SUMB_1_7_port, Y => n217);
   U355 : NAND2X1 port map( A => n1025, B => n1007, Y => n218);
   U356 : INVX2 port map( A => n218, Y => ab_3_8_port);
   U357 : XOR2X1 port map( A => n269, B => n219, Y => SUMB_3_12_port);
   U358 : XNOR2X1 port map( A => CARRYB_2_12_port, B => ab_3_12_port, Y => n219
                           );
   U359 : INVX2 port map( A => CARRYB_8_9_port, Y => n220);
   U360 : AND2X2 port map( A => n148, B => ab_1_11_port, Y => n222);
   U361 : XOR2X1 port map( A => n615, B => SUMB_2_9_port, Y => SUMB_3_8_port);
   U362 : BUFX2 port map( A => n895, Y => n225);
   U363 : XOR2X1 port map( A => n226, B => SUMB_6_8_port, Y => SUMB_7_7_port);
   U364 : XNOR2X1 port map( A => CARRYB_6_7_port, B => n440, Y => n226);
   U365 : INVX1 port map( A => SUMB_15_5_port, Y => n227);
   U366 : INVX1 port map( A => n227, Y => n228);
   U367 : XNOR2X1 port map( A => n229, B => n214, Y => SUMB_4_11_port);
   U368 : XNOR2X1 port map( A => CARRYB_3_11_port, B => ab_4_11_port, Y => n229
                           );
   U369 : INVX1 port map( A => n445, Y => n230);
   U370 : NAND3X1 port map( A => n576, B => n578, C => n577, Y => n231);
   U371 : XNOR2X1 port map( A => n232, B => SUMB_2_12_port, Y => SUMB_3_11_port
                           );
   U372 : XNOR2X1 port map( A => CARRYB_2_11_port, B => ab_3_11_port, Y => n232
                           );
   U373 : XOR2X1 port map( A => n975, B => ab_2_12_port, Y => n252);
   U374 : INVX1 port map( A => n975, Y => CARRYB_1_12_port);
   U375 : XOR2X1 port map( A => CARRYB_5_4_port, B => ab_6_4_port, Y => n233);
   U376 : XNOR2X1 port map( A => n234, B => n96, Y => SUMB_4_5_port);
   U377 : BUFX2 port map( A => n601, Y => n237);
   U378 : NAND3X1 port map( A => n872, B => n873, C => n874, Y => n238);
   U379 : INVX1 port map( A => n1006, Y => n239);
   U380 : BUFX2 port map( A => CARRYB_10_0_port, Y => n240);
   U381 : BUFX2 port map( A => n663, Y => n241);
   U382 : INVX1 port map( A => n486, Y => n242);
   U383 : INVX1 port map( A => n242, Y => n243);
   U384 : NAND3X1 port map( A => n822, B => n823, C => n824, Y => n245);
   U385 : NAND3X1 port map( A => n828, B => n830, C => n829, Y => n246);
   U386 : XOR2X1 port map( A => n411, B => n412, Y => n247);
   U387 : AND2X2 port map( A => B(15), B => n1020, Y => ab_0_15_port);
   U388 : XOR2X1 port map( A => CARRYB_6_10_port, B => n248, Y => n750);
   U389 : INVX2 port map( A => SUMB_9_8_port, Y => n736);
   U390 : XOR2X1 port map( A => n249, B => n250, Y => SUMB_6_11_port);
   U391 : XNOR2X1 port map( A => ab_6_11_port, B => CARRYB_5_11_port, Y => n249
                           );
   U392 : INVX2 port map( A => SUMB_5_12_port, Y => n250);
   U393 : XNOR2X1 port map( A => n252, B => SUMB_1_13_port, Y => SUMB_2_12_port
                           );
   U394 : NAND2X1 port map( A => ab_8_6_port, B => CARRYB_7_6_port, Y => n254);
   U395 : NAND2X1 port map( A => SUMB_7_7_port, B => ab_8_6_port, Y => n255);
   U396 : NAND2X1 port map( A => CARRYB_7_6_port, B => SUMB_7_7_port, Y => n256
                           );
   U397 : NAND3X1 port map( A => n254, B => n255, C => n256, Y => 
                           CARRYB_8_6_port);
   U398 : NAND2X1 port map( A => n204, B => ab_9_5_port, Y => n257);
   U399 : NAND2X1 port map( A => SUMB_8_6_port, B => ab_9_5_port, Y => n258);
   U400 : NAND2X1 port map( A => n204, B => SUMB_8_6_port, Y => n259);
   U401 : NAND3X1 port map( A => n257, B => n258, C => n259, Y => 
                           CARRYB_9_5_port);
   U402 : NAND3X1 port map( A => n641, B => n642, C => n643, Y => n260);
   U403 : XOR2X1 port map( A => CARRYB_4_7_port, B => n261, Y => n543);
   U404 : NAND2X1 port map( A => ab_6_5_port, B => n263, Y => n264);
   U405 : NAND2X1 port map( A => n262, B => n245, Y => n265);
   U406 : NAND2X1 port map( A => n264, B => n265, Y => n700);
   U407 : INVX1 port map( A => ab_6_5_port, Y => n262);
   U408 : INVX1 port map( A => CARRYB_5_5_port, Y => n263);
   U409 : INVX4 port map( A => B(12), Y => n1014);
   U410 : INVX2 port map( A => CARRYB_5_7_port, Y => n272);
   U411 : BUFX4 port map( A => A(0), Y => n266);
   U412 : INVX2 port map( A => A(0), Y => n1020);
   U413 : XNOR2X1 port map( A => n267, B => n268, Y => SUMB_14_3_port);
   U414 : INVX2 port map( A => SUMB_13_4_port, Y => n268);
   U415 : INVX2 port map( A => SUMB_2_13_port, Y => n269);
   U416 : NAND3X1 port map( A => n843, B => n845, C => n844, Y => n270);
   U417 : XNOR2X1 port map( A => n273, B => n274, Y => SUMB_13_3_port);
   U418 : XOR2X1 port map( A => CARRYB_12_3_port, B => ab_13_3_port, Y => n273)
                           ;
   U419 : XNOR2X1 port map( A => n339, B => n414, Y => n274);
   U420 : INVX1 port map( A => SUMB_7_2_port, Y => n373);
   U421 : NAND3X1 port map( A => n661, B => n662, C => n241, Y => n275);
   U422 : NAND3X1 port map( A => n717, B => n718, C => n719, Y => n276);
   U423 : NAND3X1 port map( A => n602, B => n603, C => n604, Y => n277);
   U424 : NAND3X1 port map( A => n878, B => n879, C => n880, Y => n278);
   U425 : NAND3X1 port map( A => n537, B => n536, C => n538, Y => n279);
   U426 : BUFX2 port map( A => n793, Y => n280);
   U427 : XNOR2X1 port map( A => n281, B => SUMB_11_8_port, Y => SUMB_12_7_port
                           );
   U428 : XNOR2X1 port map( A => CARRYB_11_7_port, B => ab_12_7_port, Y => n281
                           );
   U429 : XOR2X1 port map( A => ab_14_7_port, B => CARRYB_13_7_port, Y => n282)
                           ;
   U430 : XOR2X1 port map( A => n282, B => SUMB_13_8_port, Y => SUMB_14_7_port)
                           ;
   U431 : XOR2X1 port map( A => ab_15_6_port, B => CARRYB_14_6_port, Y => n283)
                           ;
   U432 : XOR2X1 port map( A => n283, B => SUMB_14_7_port, Y => SUMB_15_6_port)
                           ;
   U433 : NAND2X1 port map( A => ab_14_7_port, B => CARRYB_13_7_port, Y => n284
                           );
   U434 : NAND2X1 port map( A => ab_14_7_port, B => SUMB_13_8_port, Y => n285);
   U435 : NAND2X1 port map( A => CARRYB_13_7_port, B => SUMB_13_8_port, Y => 
                           n286);
   U436 : NAND3X1 port map( A => n284, B => n285, C => n286, Y => 
                           CARRYB_14_7_port);
   U437 : NAND2X1 port map( A => ab_15_6_port, B => CARRYB_14_6_port, Y => n287
                           );
   U438 : NAND2X1 port map( A => ab_15_6_port, B => SUMB_14_7_port, Y => n288);
   U439 : NAND2X1 port map( A => CARRYB_14_6_port, B => SUMB_14_7_port, Y => 
                           n289);
   U440 : NAND3X1 port map( A => n287, B => n288, C => n289, Y => 
                           CARRYB_15_6_port);
   U441 : XOR2X1 port map( A => CARRYB_11_8_port, B => ab_12_8_port, Y => n290)
                           ;
   U442 : XOR2X1 port map( A => SUMB_11_9_port, B => n290, Y => SUMB_12_8_port)
                           ;
   U443 : NAND2X1 port map( A => SUMB_11_9_port, B => n213, Y => n291);
   U444 : NAND2X1 port map( A => SUMB_11_9_port, B => ab_12_8_port, Y => n292);
   U445 : NAND2X1 port map( A => n213, B => ab_12_8_port, Y => n293);
   U446 : NAND3X1 port map( A => n292, B => n291, C => n293, Y => 
                           CARRYB_12_8_port);
   U447 : BUFX2 port map( A => CARRYB_4_12_port, Y => n294);
   U448 : NAND3X1 port map( A => n684, B => n685, C => n686, Y => n295);
   U449 : INVX2 port map( A => SUMB_1_10_port, Y => n337);
   U450 : XOR2X1 port map( A => CARRYB_13_5_port, B => ab_14_5_port, Y => n332)
                           ;
   U451 : XNOR2X1 port map( A => n296, B => n736, Y => SUMB_10_7_port);
   U452 : XOR2X1 port map( A => CARRYB_9_7_port, B => ab_10_7_port, Y => n296);
   U453 : XNOR2X1 port map( A => CARRYB_10_5_port, B => n298, Y => n598);
   U454 : NAND3X1 port map( A => n893, B => n225, C => n187, Y => n299);
   U455 : XNOR2X1 port map( A => n726, B => n300, Y => SUMB_6_9_port);
   U456 : INVX8 port map( A => B(15), Y => n1049);
   U457 : XOR2X1 port map( A => CARRYB_10_4_port, B => n301, Y => n312);
   U458 : NAND3X1 port map( A => n825, B => n826, C => n827, Y => n302);
   U459 : NAND3X1 port map( A => n832, B => n831, C => n833, Y => n303);
   U460 : XOR2X1 port map( A => SUMB_4_13_port, B => ab_5_12_port, Y => n304);
   U461 : XOR2X1 port map( A => n304, B => n294, Y => SUMB_5_12_port);
   U462 : NAND2X1 port map( A => CARRYB_4_12_port, B => SUMB_4_13_port, Y => 
                           n305);
   U463 : NAND2X1 port map( A => CARRYB_4_12_port, B => ab_5_12_port, Y => n306
                           );
   U464 : NAND2X1 port map( A => SUMB_4_13_port, B => ab_5_12_port, Y => n307);
   U465 : NAND3X1 port map( A => n307, B => n305, C => n306, Y => 
                           CARRYB_5_12_port);
   U466 : NAND2X1 port map( A => SUMB_1_14_port, B => CARRYB_1_13_port, Y => 
                           n308);
   U467 : NAND2X1 port map( A => CARRYB_1_13_port, B => ab_2_13_port, Y => n309
                           );
   U468 : NAND2X1 port map( A => n151, B => ab_2_13_port, Y => n310);
   U469 : NAND3X1 port map( A => n309, B => n308, C => n310, Y => 
                           CARRYB_2_13_port);
   U470 : NAND3X1 port map( A => n804, B => n805, C => n806, Y => n313);
   U471 : INVX2 port map( A => n1021, Y => n846);
   U472 : NAND2X1 port map( A => ab_0_8_port, B => n439, Y => n314);
   U473 : BUFX2 port map( A => SUMB_15_0_port, Y => n315);
   U474 : NAND3X1 port map( A => n500, B => n501, C => n502, Y => n316);
   U475 : XOR2X1 port map( A => SUMB_15_6_port, B => n317, Y => A1_19_port);
   U476 : XNOR2X1 port map( A => n319, B => SUMB_7_12_port, Y => SUMB_8_11_port
                           );
   U477 : XNOR2X1 port map( A => ab_8_11_port, B => CARRYB_7_11_port, Y => n319
                           );
   U478 : XOR2X1 port map( A => n474, B => n320, Y => SUMB_13_1_port);
   U479 : BUFX2 port map( A => A(1), Y => n322);
   U480 : INVX1 port map( A => A(1), Y => n1021);
   U481 : XNOR2X1 port map( A => ab_7_12_port, B => n712, Y => n680);
   U482 : INVX1 port map( A => n712, Y => n713);
   U483 : INVX1 port map( A => n441, Y => n442);
   U484 : XNOR2X1 port map( A => n323, B => n77, Y => SUMB_2_10_port);
   U485 : XNOR2X1 port map( A => SUMB_1_11_port, B => ab_2_10_port, Y => n323);
   U486 : XNOR2X1 port map( A => n324, B => CARRYB_12_8_port, Y => n457);
   U487 : XNOR2X1 port map( A => n325, B => n326, Y => SUMB_12_2_port);
   U488 : XOR2X1 port map( A => CARRYB_11_2_port, B => ab_12_2_port, Y => n325)
                           ;
   U489 : XNOR2X1 port map( A => n10, B => n374, Y => n326);
   U490 : XNOR2X1 port map( A => n327, B => SUMB_2_14_port, Y => SUMB_3_13_port
                           );
   U491 : XNOR2X1 port map( A => ab_3_13_port, B => CARRYB_2_13_port, Y => n327
                           );
   U492 : NAND3X1 port map( A => n599, B => n600, C => n237, Y => n328);
   U493 : NAND3X1 port map( A => n896, B => n897, C => n24, Y => n329);
   U494 : NAND3X1 port map( A => n658, B => n660, C => n659, Y => n330);
   U495 : XOR2X1 port map( A => n763, B => n374, Y => n331);
   U496 : XOR2X1 port map( A => n332, B => SUMB_13_6_port, Y => SUMB_14_5_port)
                           ;
   U497 : NAND2X1 port map( A => SUMB_13_6_port, B => n99, Y => n333);
   U498 : NAND2X1 port map( A => SUMB_13_6_port, B => ab_14_5_port, Y => n334);
   U499 : NAND2X1 port map( A => n99, B => ab_14_5_port, Y => n335);
   U500 : NAND3X1 port map( A => n334, B => n333, C => n335, Y => 
                           CARRYB_14_5_port);
   U501 : NAND3X1 port map( A => n891, B => n890, C => n892, Y => n336);
   U502 : XOR2X1 port map( A => n338, B => n337, Y => SUMB_2_9_port);
   U503 : XOR2X1 port map( A => n974, B => ab_2_9_port, Y => n338);
   U504 : XOR2X1 port map( A => CARRYB_10_3_port, B => ab_11_3_port, Y => n763)
                           ;
   U505 : XOR2X1 port map( A => n339, B => n414, Y => SUMB_12_4_port);
   U506 : XOR2X1 port map( A => SUMB_1_3_port, B => ab_2_2_port, Y => n340);
   U507 : XOR2X1 port map( A => n63, B => n340, Y => SUMB_2_2_port);
   U508 : NAND2X1 port map( A => n63, B => SUMB_1_3_port, Y => n341);
   U509 : NAND2X1 port map( A => n63, B => ab_2_2_port, Y => n342);
   U510 : NAND2X1 port map( A => SUMB_1_3_port, B => ab_2_2_port, Y => n343);
   U511 : NAND3X1 port map( A => n342, B => n341, C => n343, Y => 
                           CARRYB_2_2_port);
   U512 : NAND3X1 port map( A => n851, B => n850, C => n852, Y => n344);
   U513 : BUFX2 port map( A => CARRYB_13_0_port, Y => n345);
   U514 : XNOR2X1 port map( A => n346, B => n347, Y => SUMB_5_5_port);
   U515 : XOR2X1 port map( A => CARRYB_4_5_port, B => ab_5_5_port, Y => n346);
   U516 : INVX2 port map( A => SUMB_4_6_port, Y => n347);
   U517 : NAND3X1 port map( A => n875, B => n876, C => n877, Y => n348);
   U518 : NAND3X1 port map( A => n744, B => n745, C => n746, Y => n349);
   U519 : INVX2 port map( A => SUMB_11_5_port, Y => n414);
   U520 : XOR2X1 port map( A => ab_3_14_port, B => ab_2_15_port, Y => n350);
   U521 : XOR2X1 port map( A => n350, B => CARRYB_2_14_port, Y => 
                           SUMB_3_14_port);
   U522 : NAND2X1 port map( A => CARRYB_2_14_port, B => ab_3_14_port, Y => n351
                           );
   U523 : NAND2X1 port map( A => CARRYB_2_14_port, B => ab_2_15_port, Y => n352
                           );
   U524 : NAND2X1 port map( A => ab_3_14_port, B => ab_2_15_port, Y => n353);
   U525 : NAND3X1 port map( A => n352, B => n351, C => n353, Y => 
                           CARRYB_3_14_port);
   U526 : XOR2X1 port map( A => CARRYB_14_7_port, B => ab_15_7_port, Y => n354)
                           ;
   U527 : XOR2X1 port map( A => SUMB_14_8_port, B => n354, Y => SUMB_15_7_port)
                           ;
   U528 : NAND2X1 port map( A => SUMB_14_8_port, B => CARRYB_14_7_port, Y => 
                           n355);
   U529 : NAND2X1 port map( A => SUMB_14_8_port, B => ab_15_7_port, Y => n356);
   U530 : NAND2X1 port map( A => CARRYB_14_7_port, B => ab_15_7_port, Y => n357
                           );
   U531 : NAND3X1 port map( A => n356, B => n355, C => n357, Y => 
                           CARRYB_15_7_port);
   U532 : XOR2X1 port map( A => CARRYB_11_10_port, B => ab_12_10_port, Y => 
                           n358);
   U533 : XOR2X1 port map( A => SUMB_11_11_port, B => n358, Y => 
                           SUMB_12_10_port);
   U534 : NAND2X1 port map( A => SUMB_11_11_port, B => CARRYB_11_10_port, Y => 
                           n359);
   U535 : NAND2X1 port map( A => SUMB_11_11_port, B => ab_12_10_port, Y => n360
                           );
   U536 : NAND2X1 port map( A => CARRYB_11_10_port, B => ab_12_10_port, Y => 
                           n361);
   U537 : NAND3X1 port map( A => n360, B => n359, C => n361, Y => 
                           CARRYB_12_10_port);
   U538 : XOR2X1 port map( A => ab_8_13_port, B => CARRYB_7_13_port, Y => n362)
                           ;
   U539 : XOR2X1 port map( A => n362, B => SUMB_7_14_port, Y => SUMB_8_13_port)
                           ;
   U540 : NAND2X1 port map( A => ab_8_13_port, B => CARRYB_7_13_port, Y => n363
                           );
   U541 : NAND2X1 port map( A => ab_8_13_port, B => SUMB_7_14_port, Y => n364);
   U542 : NAND2X1 port map( A => CARRYB_7_13_port, B => SUMB_7_14_port, Y => 
                           n365);
   U543 : NAND3X1 port map( A => n363, B => n364, C => n365, Y => 
                           CARRYB_8_13_port);
   U544 : XOR2X1 port map( A => ab_9_13_port, B => SUMB_8_14_port, Y => n366);
   U545 : XOR2X1 port map( A => n366, B => CARRYB_8_13_port, Y => 
                           SUMB_9_13_port);
   U546 : NAND2X1 port map( A => ab_9_13_port, B => SUMB_8_14_port, Y => n367);
   U547 : NAND2X1 port map( A => ab_9_13_port, B => CARRYB_8_13_port, Y => n368
                           );
   U548 : NAND2X1 port map( A => SUMB_8_14_port, B => CARRYB_8_13_port, Y => 
                           n369);
   U549 : NAND3X1 port map( A => n367, B => n368, C => n369, Y => 
                           CARRYB_9_13_port);
   U550 : BUFX2 port map( A => n36, Y => n370);
   U551 : NAND3X1 port map( A => n753, B => n754, C => n752, Y => n371);
   U552 : XNOR2X1 port map( A => n372, B => SUMB_4_4_port, Y => SUMB_5_3_port);
   U553 : XOR2X1 port map( A => n949, B => ab_5_3_port, Y => n372);
   U554 : XNOR2X1 port map( A => n931, B => n373, Y => SUMB_8_1_port);
   U555 : XOR2X1 port map( A => n376, B => n426, Y => n374);
   U556 : INVX1 port map( A => SUMB_7_4_port, Y => n375);
   U557 : XOR2X1 port map( A => n376, B => n426, Y => SUMB_10_4_port);
   U558 : AND2X2 port map( A => n846, B => B(1), Y => ab_1_1_port);
   U559 : XNOR2X1 port map( A => n449, B => n377, Y => SUMB_10_3_port);
   U560 : INVX2 port map( A => SUMB_9_4_port, Y => n377);
   U561 : NAND2X1 port map( A => n528, B => n78, Y => n977);
   U562 : NAND3X1 port map( A => n814, B => n813, C => n815, Y => n378);
   U563 : NAND3X1 port map( A => n607, B => n605, C => n11, Y => n379);
   U564 : NAND3X1 port map( A => n781, B => n782, C => n783, Y => n380);
   U565 : NAND3X1 port map( A => n881, B => n33, C => n882, Y => n381);
   U566 : INVX1 port map( A => CARRYB_2_10_port, Y => n909);
   U567 : NAND2X1 port map( A => SUMB_10_5_port, B => n203, Y => n382);
   U568 : NAND2X1 port map( A => SUMB_10_5_port, B => ab_11_4_port, Y => n383);
   U569 : NAND2X1 port map( A => n203, B => ab_11_4_port, Y => n384);
   U570 : NAND3X1 port map( A => n384, B => n382, C => n383, Y => 
                           CARRYB_11_4_port);
   U571 : NAND3X1 port map( A => n899, B => n900, C => n901, Y => n385);
   U572 : NAND3X1 port map( A => n747, B => n119, C => n749, Y => n386);
   U573 : NAND3X1 port map( A => n590, B => n591, C => n592, Y => n387);
   U574 : NAND3X1 port map( A => n784, B => n785, C => n786, Y => n388);
   U575 : INVX1 port map( A => SUMB_13_3_port, Y => n425);
   U576 : XOR2X1 port map( A => CARRYB_10_8_port, B => ab_11_8_port, Y => n389)
                           ;
   U577 : XOR2X1 port map( A => SUMB_10_9_port, B => n389, Y => SUMB_11_8_port)
                           ;
   U578 : NAND2X1 port map( A => SUMB_10_9_port, B => CARRYB_10_8_port, Y => 
                           n390);
   U579 : NAND2X1 port map( A => SUMB_10_9_port, B => ab_11_8_port, Y => n391);
   U580 : NAND2X1 port map( A => CARRYB_10_8_port, B => ab_11_8_port, Y => n392
                           );
   U581 : NAND3X1 port map( A => n391, B => n390, C => n392, Y => 
                           CARRYB_11_8_port);
   U582 : NAND3X1 port map( A => n697, B => n699, C => n123, Y => n393);
   U583 : NAND3X1 port map( A => n652, B => n653, C => n654, Y => n394);
   U584 : XNOR2X1 port map( A => n648, B => n395, Y => SUMB_3_4_port);
   U585 : INVX1 port map( A => SUMB_2_5_port, Y => n395);
   U586 : BUFX2 port map( A => n1025, Y => n396);
   U587 : XOR2X1 port map( A => CARRYB_3_3_port, B => ab_4_3_port, Y => n397);
   U588 : XOR2X1 port map( A => SUMB_3_4_port, B => n397, Y => SUMB_4_3_port);
   U589 : NAND2X1 port map( A => SUMB_3_4_port, B => CARRYB_3_3_port, Y => n398
                           );
   U590 : NAND2X1 port map( A => SUMB_3_4_port, B => ab_4_3_port, Y => n399);
   U591 : NAND2X1 port map( A => CARRYB_3_3_port, B => ab_4_3_port, Y => n400);
   U592 : NAND3X1 port map( A => n400, B => n399, C => n398, Y => 
                           CARRYB_4_3_port);
   U593 : INVX1 port map( A => CARRYB_4_3_port, Y => n949);
   U594 : INVX4 port map( A => A(3), Y => n1024);
   U595 : AND2X2 port map( A => n236, B => B(7), Y => n435);
   U596 : XOR2X1 port map( A => SUMB_3_10_port, B => n401, Y => n454);
   U597 : XOR2X1 port map( A => n174, B => ab_10_2_port, Y => n402);
   U598 : XOR2X1 port map( A => SUMB_9_3_port, B => n402, Y => SUMB_10_2_port);
   U599 : NAND2X1 port map( A => SUMB_9_3_port, B => CARRYB_9_2_port, Y => n403
                           );
   U600 : NAND2X1 port map( A => SUMB_9_3_port, B => ab_10_2_port, Y => n404);
   U601 : NAND2X1 port map( A => CARRYB_9_2_port, B => ab_10_2_port, Y => n405)
                           ;
   U602 : NAND3X1 port map( A => n404, B => n403, C => n405, Y => 
                           CARRYB_10_2_port);
   U603 : XNOR2X1 port map( A => ab_1_5_port, B => n406, Y => SUMB_1_5_port);
   U604 : NAND2X1 port map( A => B(6), B => n987, Y => n406);
   U605 : NAND2X1 port map( A => SUMB_4_12_port, B => n16, Y => n407);
   U606 : NAND2X1 port map( A => SUMB_4_12_port, B => ab_5_11_port, Y => n408);
   U607 : NAND2X1 port map( A => n16, B => ab_5_11_port, Y => n409);
   U608 : NAND3X1 port map( A => n408, B => n407, C => n409, Y => 
                           CARRYB_5_11_port);
   U609 : INVX2 port map( A => CARRYB_5_6_port, Y => n445);
   U610 : XOR2X1 port map( A => n410, B => n534, Y => SUMB_8_4_port);
   U611 : INVX1 port map( A => SUMB_3_9_port, Y => n411);
   U612 : XNOR2X1 port map( A => CARRYB_3_8_port, B => ab_4_8_port, Y => n412);
   U613 : NAND3X1 port map( A => n453, B => n452, C => n451, Y => n413);
   U614 : BUFX2 port map( A => n75, Y => n415);
   U615 : XOR2X1 port map( A => ab_8_12_port, B => CARRYB_7_12_port, Y => n416)
                           ;
   U616 : XOR2X1 port map( A => n416, B => SUMB_7_13_port, Y => SUMB_8_12_port)
                           ;
   U617 : XOR2X1 port map( A => ab_9_11_port, B => CARRYB_8_11_port, Y => n417)
                           ;
   U618 : XOR2X1 port map( A => n417, B => SUMB_8_12_port, Y => SUMB_9_11_port)
                           ;
   U619 : NAND2X1 port map( A => ab_8_12_port, B => CARRYB_7_12_port, Y => n418
                           );
   U620 : NAND2X1 port map( A => ab_8_12_port, B => SUMB_7_13_port, Y => n419);
   U621 : NAND2X1 port map( A => CARRYB_7_12_port, B => SUMB_7_13_port, Y => 
                           n420);
   U622 : NAND3X1 port map( A => n418, B => n419, C => n420, Y => 
                           CARRYB_8_12_port);
   U623 : NAND2X1 port map( A => ab_9_11_port, B => n295, Y => n421);
   U624 : NAND2X1 port map( A => ab_9_11_port, B => SUMB_8_12_port, Y => n422);
   U625 : NAND2X1 port map( A => n295, B => SUMB_8_12_port, Y => n423);
   U626 : NAND3X1 port map( A => n421, B => n422, C => n423, Y => 
                           CARRYB_9_11_port);
   U627 : INVX2 port map( A => n986, Y => n511);
   U628 : XOR2X1 port map( A => SUMB_12_7_port, B => n424, Y => SUMB_13_6_port)
                           ;
   U629 : XOR2X1 port map( A => n575, B => n425, Y => SUMB_14_2_port);
   U630 : INVX2 port map( A => SUMB_9_5_port, Y => n426);
   U631 : XOR2X1 port map( A => CARRYB_14_3_port, B => ab_15_3_port, Y => n427)
                           ;
   U632 : XOR2X1 port map( A => SUMB_14_4_port, B => n427, Y => SUMB_15_3_port)
                           ;
   U633 : NAND2X1 port map( A => SUMB_14_4_port, B => n275, Y => n428);
   U634 : NAND2X1 port map( A => SUMB_14_4_port, B => ab_15_3_port, Y => n429);
   U635 : NAND2X1 port map( A => n275, B => ab_15_3_port, Y => n430);
   U636 : NAND3X1 port map( A => n429, B => n428, C => n430, Y => 
                           CARRYB_15_3_port);
   U637 : INVX1 port map( A => B(7), Y => n1004);
   U638 : BUFX2 port map( A => SUMB_10_1_port, Y => n432);
   U639 : NAND3X1 port map( A => n630, B => n629, C => n631, Y => n433);
   U640 : XNOR2X1 port map( A => SUMB_4_3_port, B => n434, Y => SUMB_5_2_port);
   U641 : XNOR2X1 port map( A => CARRYB_4_2_port, B => ab_5_2_port, Y => n434);
   U642 : NAND2X1 port map( A => ab_3_8_port, B => n436, Y => n437);
   U643 : NAND2X1 port map( A => n218, B => n126, Y => n438);
   U644 : NAND2X1 port map( A => n437, B => n438, Y => n615);
   U645 : AND2X2 port map( A => B(7), B => n511, Y => n439);
   U646 : BUFX2 port map( A => SUMB_12_1_port, Y => n443);
   U647 : NAND2X1 port map( A => n445, B => ab_6_6_port, Y => n446);
   U648 : NAND2X1 port map( A => n444, B => n193, Y => n447);
   U649 : NAND2X1 port map( A => n446, B => n447, Y => n923);
   U650 : INVX1 port map( A => ab_6_6_port, Y => n444);
   U651 : XNOR2X1 port map( A => ab_8_5_port, B => CARRYB_7_5_port, Y => n448);
   U652 : XOR2X1 port map( A => SUMB_5_4_port, B => ab_6_3_port, Y => n450);
   U653 : XOR2X1 port map( A => n15, B => n450, Y => SUMB_6_3_port);
   U654 : NAND2X1 port map( A => SUMB_5_4_port, B => CARRYB_5_3_port, Y => n451
                           );
   U655 : NAND2X1 port map( A => CARRYB_5_3_port, B => ab_6_3_port, Y => n452);
   U656 : NAND2X1 port map( A => SUMB_5_4_port, B => ab_6_3_port, Y => n453);
   U657 : NAND3X1 port map( A => n453, B => n451, C => n452, Y => 
                           CARRYB_6_3_port);
   U658 : XNOR2X1 port map( A => n454, B => n978, Y => SUMB_4_9_port);
   U659 : XOR2X1 port map( A => n455, B => n608, Y => SUMB_9_2_port);
   U660 : XNOR2X1 port map( A => ab_9_2_port, B => n197, Y => n455);
   U661 : XOR2X1 port map( A => ab_12_9_port, B => CARRYB_11_9_port, Y => n456)
                           ;
   U662 : XOR2X1 port map( A => n456, B => SUMB_11_10_port, Y => SUMB_12_9_port
                           );
   U663 : XOR2X1 port map( A => n457, B => SUMB_12_9_port, Y => SUMB_13_8_port)
                           ;
   U664 : NAND2X1 port map( A => ab_12_9_port, B => CARRYB_11_9_port, Y => n458
                           );
   U665 : NAND2X1 port map( A => ab_12_9_port, B => SUMB_11_10_port, Y => n459)
                           ;
   U666 : NAND2X1 port map( A => CARRYB_11_9_port, B => SUMB_11_10_port, Y => 
                           n460);
   U667 : NAND3X1 port map( A => n458, B => n459, C => n460, Y => 
                           CARRYB_12_9_port);
   U668 : NAND2X1 port map( A => ab_13_8_port, B => CARRYB_12_8_port, Y => n461
                           );
   U669 : NAND2X1 port map( A => ab_13_8_port, B => SUMB_12_9_port, Y => n462);
   U670 : NAND2X1 port map( A => CARRYB_12_8_port, B => SUMB_12_9_port, Y => 
                           n463);
   U671 : NAND3X1 port map( A => n461, B => n462, C => n463, Y => 
                           CARRYB_13_8_port);
   U672 : XNOR2X1 port map( A => ab_0_9_port, B => n464, Y => SUMB_1_8_port);
   U673 : NAND2X1 port map( A => n1007, B => n514, Y => n464);
   U674 : NAND2X1 port map( A => ab_9_9_port, B => n221, Y => n465);
   U675 : NAND2X1 port map( A => SUMB_8_10_port, B => ab_9_9_port, Y => n466);
   U676 : NAND2X1 port map( A => n221, B => SUMB_8_10_port, Y => n467);
   U677 : NAND3X1 port map( A => n465, B => n466, C => n467, Y => 
                           CARRYB_9_9_port);
   U678 : NAND2X1 port map( A => ab_10_8_port, B => n349, Y => n468);
   U679 : NAND2X1 port map( A => ab_10_8_port, B => SUMB_9_9_port, Y => n469);
   U680 : NAND2X1 port map( A => n349, B => SUMB_9_9_port, Y => n470);
   U681 : NAND3X1 port map( A => n468, B => n469, C => n470, Y => 
                           CARRYB_10_8_port);
   U682 : INVX1 port map( A => n1017, Y => n1038);
   U683 : XNOR2X1 port map( A => n471, B => SUMB_3_13_port, Y => SUMB_4_12_port
                           );
   U684 : XOR2X1 port map( A => ab_4_12_port, B => n593, Y => n471);
   U685 : NAND2X1 port map( A => n487, B => n485, Y => n472);
   U686 : NAND2X1 port map( A => n243, B => n473, Y => n980);
   U687 : INVX4 port map( A => B(13), Y => n1016);
   U688 : XNOR2X1 port map( A => n371, B => ab_13_1_port, Y => n474);
   U689 : NAND3X1 port map( A => n12, B => n88, C => n637, Y => n475);
   U690 : BUFX2 port map( A => CARRYB_4_6_port, Y => n476);
   U691 : INVX4 port map( A => B(11), Y => n1012);
   U692 : XOR2X1 port map( A => SUMB_4_7_port, B => ab_5_6_port, Y => n477);
   U693 : XOR2X1 port map( A => n477, B => n476, Y => SUMB_5_6_port);
   U694 : NAND2X1 port map( A => SUMB_4_7_port, B => CARRYB_4_6_port, Y => n478
                           );
   U695 : NAND2X1 port map( A => CARRYB_4_6_port, B => ab_5_6_port, Y => n479);
   U696 : NAND2X1 port map( A => ab_5_6_port, B => SUMB_4_7_port, Y => n480);
   U697 : NAND3X1 port map( A => n478, B => n479, C => n480, Y => 
                           CARRYB_5_6_port);
   U698 : NAND2X1 port map( A => SUMB_14_1_port, B => n316, Y => n481);
   U699 : NAND2X1 port map( A => SUMB_14_1_port, B => ab_15_0_port, Y => n482);
   U700 : NAND2X1 port map( A => n316, B => ab_15_0_port, Y => n483);
   U701 : NAND3X1 port map( A => n483, B => n481, C => n482, Y => 
                           CARRYB_15_0_port);
   U702 : NAND3X1 port map( A => n914, B => n915, C => n916, Y => n484);
   U703 : NAND2X1 port map( A => n93, B => n53, Y => n485);
   U704 : NAND2X1 port map( A => n93, B => ab_12_3_port, Y => n486);
   U705 : NAND2X1 port map( A => n53, B => ab_12_3_port, Y => n487);
   U706 : NAND3X1 port map( A => n487, B => n485, C => n486, Y => 
                           CARRYB_12_3_port);
   U707 : NAND3X1 port map( A => n757, B => n756, C => n758, Y => n488);
   U708 : NAND3X1 port map( A => n623, B => n622, C => n621, Y => n489);
   U709 : NAND3X1 port map( A => n948, B => n947, C => n946, Y => n490);
   U710 : NAND3X1 port map( A => n913, B => n912, C => n911, Y => n491);
   U711 : NAND3X1 port map( A => n917, B => n918, C => n919, Y => n492);
   U712 : NAND3X1 port map( A => n579, B => n580, C => n581, Y => n493);
   U713 : NAND3X1 port map( A => n671, B => n670, C => n672, Y => n494);
   U714 : XOR2X1 port map( A => SUMB_2_2_port, B => ab_3_1_port, Y => n495);
   U715 : XOR2X1 port map( A => CARRYB_2_1_port, B => n495, Y => SUMB_3_1_port)
                           ;
   U716 : NAND2X1 port map( A => CARRYB_2_1_port, B => SUMB_2_2_port, Y => n496
                           );
   U717 : NAND2X1 port map( A => CARRYB_2_1_port, B => ab_3_1_port, Y => n497);
   U718 : NAND2X1 port map( A => SUMB_2_2_port, B => ab_3_1_port, Y => n498);
   U719 : NAND3X1 port map( A => n497, B => n496, C => n498, Y => 
                           CARRYB_3_1_port);
   U720 : XOR2X1 port map( A => n370, B => ab_14_0_port, Y => n499);
   U721 : XOR2X1 port map( A => n499, B => n345, Y => A1_12_port);
   U722 : NAND2X1 port map( A => SUMB_13_1_port, B => CARRYB_13_0_port, Y => 
                           n500);
   U723 : NAND2X1 port map( A => CARRYB_13_0_port, B => ab_14_0_port, Y => n501
                           );
   U724 : NAND2X1 port map( A => SUMB_13_1_port, B => ab_14_0_port, Y => n502);
   U725 : NAND3X1 port map( A => n501, B => n500, C => n502, Y => 
                           CARRYB_14_0_port);
   U726 : XOR2X1 port map( A => ab_2_3_port, B => SUMB_1_4_port, Y => n504);
   U727 : XOR2X1 port map( A => n970, B => n504, Y => SUMB_2_3_port);
   U728 : NAND2X1 port map( A => n970, B => ab_2_3_port, Y => n505);
   U729 : NAND2X1 port map( A => n970, B => SUMB_1_4_port, Y => n506);
   U730 : NAND2X1 port map( A => ab_2_3_port, B => SUMB_1_4_port, Y => n507);
   U731 : NAND3X1 port map( A => n506, B => n505, C => n507, Y => 
                           CARRYB_2_3_port);
   U732 : NAND2X1 port map( A => SUMB_4_3_port, B => n145, Y => n508);
   U733 : NAND2X1 port map( A => SUMB_4_3_port, B => ab_5_2_port, Y => n509);
   U734 : NAND2X1 port map( A => n145, B => ab_5_2_port, Y => n510);
   U735 : NAND3X1 port map( A => n509, B => n508, C => n510, Y => 
                           CARRYB_5_2_port);
   U736 : INVX1 port map( A => n132, Y => n1042);
   U737 : XOR2X1 port map( A => n512, B => n513, Y => SUMB_3_7_port);
   U738 : XNOR2X1 port map( A => ab_3_7_port, B => n302, Y => n512);
   U739 : INVX1 port map( A => SUMB_2_8_port, Y => n513);
   U740 : XOR2X1 port map( A => SUMB_3_2_port, B => ab_4_1_port, Y => n515);
   U741 : XOR2X1 port map( A => CARRYB_3_1_port, B => n515, Y => SUMB_4_1_port)
                           ;
   U742 : NAND2X1 port map( A => SUMB_3_2_port, B => CARRYB_3_1_port, Y => n516
                           );
   U743 : NAND2X1 port map( A => CARRYB_3_1_port, B => ab_4_1_port, Y => n517);
   U744 : NAND2X1 port map( A => SUMB_3_2_port, B => ab_4_1_port, Y => n518);
   U745 : NAND3X1 port map( A => n517, B => n516, C => n518, Y => 
                           CARRYB_4_1_port);
   U746 : XOR2X1 port map( A => n181, B => ab_2_6_port, Y => n519);
   U747 : NAND2X1 port map( A => SUMB_1_7_port, B => n181, Y => n520);
   U748 : NAND2X1 port map( A => SUMB_1_7_port, B => ab_2_6_port, Y => n521);
   U749 : NAND2X1 port map( A => n181, B => ab_2_6_port, Y => n522);
   U750 : NAND3X1 port map( A => n520, B => n521, C => n522, Y => 
                           CARRYB_2_6_port);
   U751 : NAND3X1 port map( A => n559, B => n558, C => n560, Y => n523);
   U752 : INVX1 port map( A => n1013, Y => n1040);
   U753 : AND2X2 port map( A => n999, B => n514, Y => n525);
   U754 : BUFX2 port map( A => SUMB_1_6_port, Y => n526);
   U755 : INVX1 port map( A => n1009, Y => n1041);
   U756 : NAND2X1 port map( A => SUMB_1_10_port, B => CARRYB_1_9_port, Y => 
                           n527);
   U757 : NAND2X1 port map( A => SUMB_1_10_port, B => ab_2_9_port, Y => n528);
   U758 : NAND2X1 port map( A => ab_2_9_port, B => CARRYB_1_9_port, Y => n529);
   U759 : NAND3X1 port map( A => n528, B => n527, C => n529, Y => 
                           CARRYB_2_9_port);
   U760 : XNOR2X1 port map( A => CARRYB_13_1_port, B => n530, Y => n633);
   U761 : BUFX2 port map( A => SUMB_6_3_port, Y => n531);
   U762 : XNOR2X1 port map( A => n532, B => SUMB_3_8_port, Y => SUMB_4_7_port);
   U763 : NAND3X1 port map( A => n649, B => n650, C => n651, Y => n533);
   U764 : XOR2X1 port map( A => CARRYB_10_6_port, B => ab_11_6_port, Y => n535)
                           ;
   U765 : XOR2X1 port map( A => n535, B => SUMB_10_7_port, Y => SUMB_11_6_port)
                           ;
   U766 : NAND2X1 port map( A => SUMB_10_7_port, B => n379, Y => n536);
   U767 : NAND2X1 port map( A => SUMB_10_7_port, B => ab_11_6_port, Y => n537);
   U768 : NAND2X1 port map( A => n379, B => ab_11_6_port, Y => n538);
   U769 : NAND3X1 port map( A => n537, B => n536, C => n538, Y => 
                           CARRYB_11_6_port);
   U770 : NAND3X1 port map( A => n787, B => n789, C => n788, Y => n539);
   U771 : NAND3X1 port map( A => n611, B => n610, C => n612, Y => n540);
   U772 : INVX2 port map( A => n1000, Y => n985);
   U773 : XNOR2X1 port map( A => n700, B => n541, Y => SUMB_6_5_port);
   U774 : INVX2 port map( A => SUMB_5_6_port, Y => n541);
   U775 : INVX1 port map( A => n951, Y => n939);
   U776 : INVX4 port map( A => B(9), Y => n1008);
   U777 : XNOR2X1 port map( A => n543, B => n247, Y => SUMB_5_7_port);
   U778 : NAND2X1 port map( A => ab_13_7_port, B => n19, Y => n544);
   U779 : NAND2X1 port map( A => SUMB_12_8_port, B => ab_13_7_port, Y => n545);
   U780 : NAND2X1 port map( A => n19, B => SUMB_12_8_port, Y => n546);
   U781 : NAND3X1 port map( A => n544, B => n545, C => n546, Y => 
                           CARRYB_13_7_port);
   U782 : NAND2X1 port map( A => ab_14_6_port, B => n393, Y => n547);
   U783 : NAND2X1 port map( A => SUMB_13_7_port, B => ab_14_6_port, Y => n548);
   U784 : NAND2X1 port map( A => SUMB_13_7_port, B => n393, Y => n549);
   U785 : NAND3X1 port map( A => n547, B => n548, C => n549, Y => 
                           CARRYB_14_6_port);
   U786 : NAND2X1 port map( A => SUMB_2_13_port, B => n238, Y => n550);
   U787 : NAND2X1 port map( A => SUMB_2_13_port, B => ab_3_12_port, Y => n551);
   U788 : NAND2X1 port map( A => n238, B => ab_3_12_port, Y => n552);
   U789 : NAND3X1 port map( A => n551, B => n550, C => n552, Y => 
                           CARRYB_3_12_port);
   U790 : XOR2X1 port map( A => SUMB_9_10_port, B => ab_10_9_port, Y => n553);
   U791 : XOR2X1 port map( A => n553, B => CARRYB_9_9_port, Y => SUMB_10_9_port
                           );
   U792 : NAND2X1 port map( A => CARRYB_9_9_port, B => SUMB_9_10_port, Y => 
                           n554);
   U793 : NAND2X1 port map( A => CARRYB_9_9_port, B => ab_10_9_port, Y => n555)
                           ;
   U794 : NAND2X1 port map( A => SUMB_9_10_port, B => ab_10_9_port, Y => n556);
   U795 : NAND3X1 port map( A => n555, B => n554, C => n556, Y => 
                           CARRYB_10_9_port);
   U796 : NAND3X1 port map( A => n792, B => n120, C => n280, Y => n557);
   U797 : NAND2X1 port map( A => CARRYB_3_5_port, B => SUMB_3_6_port, Y => n558
                           );
   U798 : NAND2X1 port map( A => CARRYB_3_5_port, B => ab_4_5_port, Y => n559);
   U799 : NAND2X1 port map( A => SUMB_3_6_port, B => ab_4_5_port, Y => n560);
   U800 : NAND3X1 port map( A => n560, B => n559, C => n558, Y => 
                           CARRYB_4_5_port);
   U801 : XOR2X1 port map( A => n561, B => SUMB_14_2_port, Y => SUMB_15_1_port)
                           ;
   U802 : NAND2X1 port map( A => SUMB_14_2_port, B => n475, Y => n562);
   U803 : NAND2X1 port map( A => SUMB_14_2_port, B => ab_15_1_port, Y => n563);
   U804 : NAND2X1 port map( A => n475, B => ab_15_1_port, Y => n564);
   U805 : NAND3X1 port map( A => n564, B => n562, C => n563, Y => 
                           CARRYB_15_1_port);
   U806 : NAND3X1 port map( A => n840, B => n841, C => n842, Y => n565);
   U807 : NAND3X1 port map( A => n634, B => n636, C => n635, Y => n566);
   U808 : NAND2X1 port map( A => SUMB_5_3_port, B => CARRYB_5_2_port, Y => n567
                           );
   U809 : NAND2X1 port map( A => CARRYB_5_2_port, B => ab_6_2_port, Y => n568);
   U810 : NAND2X1 port map( A => SUMB_5_3_port, B => ab_6_2_port, Y => n569);
   U811 : NAND3X1 port map( A => n568, B => n567, C => n569, Y => 
                           CARRYB_6_2_port);
   U812 : XNOR2X1 port map( A => n952, B => ab_5_1_port, Y => n857);
   U813 : INVX1 port map( A => n1015, Y => n1039);
   U814 : BUFX4 port map( A => CARRYB_3_9_port, Y => n978);
   U815 : XNOR2X1 port map( A => n570, B => SUMB_12_5_port, Y => SUMB_13_4_port
                           );
   U816 : XNOR2X1 port map( A => CARRYB_12_4_port, B => ab_13_4_port, Y => n570
                           );
   U817 : INVX1 port map( A => n593, Y => n594);
   U818 : XOR2X1 port map( A => ab_2_14_port, B => ab_1_15_port, Y => n571);
   U819 : XOR2X1 port map( A => n415, B => n571, Y => SUMB_2_14_port);
   U820 : NAND2X1 port map( A => n75, B => ab_2_14_port, Y => n572);
   U821 : NAND2X1 port map( A => n75, B => ab_1_15_port, Y => n573);
   U822 : NAND2X1 port map( A => ab_2_14_port, B => ab_1_15_port, Y => n574);
   U823 : NAND3X1 port map( A => n573, B => n572, C => n574, Y => 
                           CARRYB_2_14_port);
   U824 : XNOR2X1 port map( A => n566, B => ab_14_2_port, Y => n575);
   U825 : INVX4 port map( A => B(14), Y => n1018);
   U826 : NAND2X1 port map( A => ab_12_2_port, B => n492, Y => n576);
   U827 : NAND2X1 port map( A => n331, B => ab_12_2_port, Y => n577);
   U828 : NAND2X1 port map( A => n331, B => n492, Y => n578);
   U829 : NAND3X1 port map( A => n576, B => n578, C => n577, Y => 
                           CARRYB_12_2_port);
   U830 : NAND2X1 port map( A => ab_13_1_port, B => CARRYB_12_1_port, Y => n579
                           );
   U831 : NAND2X1 port map( A => SUMB_12_2_port, B => ab_13_1_port, Y => n580);
   U832 : NAND2X1 port map( A => SUMB_12_2_port, B => CARRYB_12_1_port, Y => 
                           n581);
   U833 : NAND3X1 port map( A => n581, B => n580, C => n579, Y => 
                           CARRYB_13_1_port);
   U834 : INVX4 port map( A => n1020, Y => n987);
   U835 : INVX1 port map( A => n909, Y => n910);
   U836 : XOR2X1 port map( A => n432, B => ab_11_0_port, Y => n582);
   U837 : XOR2X1 port map( A => n240, B => n582, Y => A1_9_port);
   U838 : NAND2X1 port map( A => CARRYB_10_0_port, B => SUMB_10_1_port, Y => 
                           n583);
   U839 : NAND2X1 port map( A => CARRYB_10_0_port, B => ab_11_0_port, Y => n584
                           );
   U840 : NAND2X1 port map( A => SUMB_10_1_port, B => ab_11_0_port, Y => n585);
   U841 : NAND3X1 port map( A => n585, B => n583, C => n584, Y => 
                           CARRYB_11_0_port);
   U842 : NAND2X1 port map( A => ab_11_7_port, B => n386, Y => n587);
   U843 : NAND2X1 port map( A => SUMB_10_8_port, B => ab_11_7_port, Y => n588);
   U844 : NAND2X1 port map( A => SUMB_10_8_port, B => n386, Y => n589);
   U845 : NAND3X1 port map( A => n587, B => n588, C => n589, Y => 
                           CARRYB_11_7_port);
   U846 : NAND2X1 port map( A => ab_12_6_port, B => n279, Y => n590);
   U847 : NAND2X1 port map( A => ab_12_6_port, B => n76, Y => n591);
   U848 : NAND2X1 port map( A => n279, B => n76, Y => n592);
   U849 : NAND3X1 port map( A => n590, B => n592, C => n591, Y => 
                           CARRYB_12_6_port);
   U850 : INVX2 port map( A => CARRYB_3_12_port, Y => n593);
   U851 : NAND2X1 port map( A => SUMB_3_9_port, B => n565, Y => n595);
   U852 : NAND2X1 port map( A => SUMB_3_9_port, B => ab_4_8_port, Y => n596);
   U853 : NAND2X1 port map( A => n565, B => ab_4_8_port, Y => n597);
   U854 : NAND3X1 port map( A => n597, B => n595, C => n596, Y => 
                           CARRYB_4_8_port);
   U855 : XOR2X1 port map( A => SUMB_10_6_port, B => n598, Y => SUMB_11_5_port)
                           ;
   U856 : NAND2X1 port map( A => ab_11_5_port, B => n276, Y => n599);
   U857 : NAND2X1 port map( A => SUMB_10_6_port, B => ab_11_5_port, Y => n600);
   U858 : NAND2X1 port map( A => SUMB_10_6_port, B => n276, Y => n601);
   U859 : NAND3X1 port map( A => n599, B => n600, C => n601, Y => 
                           CARRYB_11_5_port);
   U860 : NAND2X1 port map( A => ab_12_4_port, B => n180, Y => n602);
   U861 : NAND2X1 port map( A => ab_12_4_port, B => SUMB_11_5_port, Y => n603);
   U862 : NAND2X1 port map( A => SUMB_11_5_port, B => n180, Y => n604);
   U863 : NAND3X1 port map( A => n602, B => n603, C => n604, Y => 
                           CARRYB_12_4_port);
   U864 : NAND2X1 port map( A => SUMB_9_7_port, B => n87, Y => n605);
   U865 : NAND2X1 port map( A => SUMB_9_7_port, B => ab_10_6_port, Y => n606);
   U866 : NAND2X1 port map( A => n87, B => ab_10_6_port, Y => n607);
   U867 : NAND3X1 port map( A => n607, B => n605, C => n606, Y => 
                           CARRYB_10_6_port);
   U868 : XOR2X1 port map( A => CARRYB_11_5_port, B => ab_12_5_port, Y => n609)
                           ;
   U869 : XOR2X1 port map( A => n609, B => SUMB_11_6_port, Y => SUMB_12_5_port)
                           ;
   U870 : NAND2X1 port map( A => SUMB_11_6_port, B => n328, Y => n610);
   U871 : NAND2X1 port map( A => SUMB_11_6_port, B => ab_12_5_port, Y => n611);
   U872 : NAND2X1 port map( A => n328, B => ab_12_5_port, Y => n612);
   U873 : NAND3X1 port map( A => n612, B => n610, C => n611, Y => 
                           CARRYB_12_5_port);
   U874 : NAND3X1 port map( A => n761, B => n760, C => n762, Y => n613);
   U875 : NAND3X1 port map( A => n927, B => n928, C => n929, Y => n614);
   U876 : XOR2X1 port map( A => n443, B => ab_13_0_port, Y => n616);
   U877 : XOR2X1 port map( A => n144, B => n616, Y => A1_11_port);
   U878 : NAND2X1 port map( A => CARRYB_12_0_port, B => SUMB_12_1_port, Y => 
                           n617);
   U879 : NAND2X1 port map( A => CARRYB_12_0_port, B => ab_13_0_port, Y => n618
                           );
   U880 : NAND2X1 port map( A => SUMB_12_1_port, B => ab_13_0_port, Y => n619);
   U881 : NAND3X1 port map( A => n619, B => n617, C => n618, Y => 
                           CARRYB_13_0_port);
   U882 : NAND3X1 port map( A => n704, B => n705, C => n706, Y => n620);
   U883 : NAND2X1 port map( A => n980, B => ab_13_3_port, Y => n621);
   U884 : NAND2X1 port map( A => SUMB_12_4_port, B => ab_13_3_port, Y => n622);
   U885 : NAND2X1 port map( A => n980, B => SUMB_12_4_port, Y => n623);
   U886 : NAND3X1 port map( A => n623, B => n622, C => n621, Y => 
                           CARRYB_13_3_port);
   U887 : NAND2X1 port map( A => CARRYB_13_2_port, B => ab_14_2_port, Y => n624
                           );
   U888 : NAND2X1 port map( A => SUMB_13_3_port, B => ab_14_2_port, Y => n625);
   U889 : NAND2X1 port map( A => CARRYB_13_2_port, B => SUMB_13_3_port, Y => 
                           n626);
   U890 : NAND3X1 port map( A => n624, B => n625, C => n626, Y => 
                           CARRYB_14_2_port);
   U891 : NAND2X1 port map( A => n940, B => n941, Y => n627);
   U892 : XOR2X1 port map( A => SUMB_8_2_port, B => ab_9_1_port, Y => n628);
   U893 : XOR2X1 port map( A => n632, B => n628, Y => SUMB_9_1_port);
   U894 : NAND2X1 port map( A => SUMB_8_2_port, B => CARRYB_8_1_port, Y => n629
                           );
   U895 : NAND2X1 port map( A => CARRYB_8_1_port, B => ab_9_1_port, Y => n630);
   U896 : NAND2X1 port map( A => SUMB_8_2_port, B => ab_9_1_port, Y => n631);
   U897 : NAND3X1 port map( A => n631, B => n629, C => n630, Y => 
                           CARRYB_9_1_port);
   U898 : BUFX2 port map( A => CARRYB_8_1_port, Y => n632);
   U899 : XOR2X1 port map( A => n633, B => SUMB_13_2_port, Y => SUMB_14_1_port)
                           ;
   U900 : NAND2X1 port map( A => ab_13_2_port, B => n231, Y => n634);
   U901 : NAND2X1 port map( A => ab_13_2_port, B => SUMB_12_3_port, Y => n635);
   U902 : NAND2X1 port map( A => SUMB_12_3_port, B => n231, Y => n636);
   U903 : NAND3X1 port map( A => n634, B => n636, C => n635, Y => 
                           CARRYB_13_2_port);
   U904 : NAND2X1 port map( A => n493, B => ab_14_1_port, Y => n637);
   U905 : NAND2X1 port map( A => SUMB_13_2_port, B => ab_14_1_port, Y => n638);
   U906 : NAND2X1 port map( A => SUMB_13_2_port, B => n493, Y => n639);
   U907 : NAND3X1 port map( A => n637, B => n639, C => n638, Y => 
                           CARRYB_14_1_port);
   U908 : NOR2X1 port map( A => n1022, B => n998, Y => ab_2_4_port);
   U909 : XOR2X1 port map( A => ab_4_4_port, B => n394, Y => n640);
   U910 : XOR2X1 port map( A => n640, B => n196, Y => SUMB_4_4_port);
   U911 : NAND2X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, Y => n641);
   U912 : NAND2X1 port map( A => ab_4_4_port, B => SUMB_3_5_port, Y => n642);
   U913 : NAND2X1 port map( A => CARRYB_3_4_port, B => SUMB_3_5_port, Y => n643
                           );
   U914 : NAND2X1 port map( A => ab_5_3_port, B => n185, Y => n644);
   U915 : NAND2X1 port map( A => SUMB_4_4_port, B => ab_5_3_port, Y => n645);
   U916 : NAND2X1 port map( A => n185, B => SUMB_4_4_port, Y => n646);
   U917 : NAND3X1 port map( A => n645, B => n644, C => n646, Y => 
                           CARRYB_5_3_port);
   U918 : XOR2X1 port map( A => n62, B => n950, Y => n647);
   U919 : XOR2X1 port map( A => n647, B => n526, Y => SUMB_2_5_port);
   U920 : XOR2X1 port map( A => CARRYB_2_4_port, B => ab_3_4_port, Y => n648);
   U921 : NAND2X1 port map( A => n62, B => n950, Y => n649);
   U922 : NAND2X1 port map( A => SUMB_1_6_port, B => n62, Y => n650);
   U923 : NAND2X1 port map( A => n950, B => SUMB_1_6_port, Y => n651);
   U924 : NAND3X1 port map( A => n649, B => n650, C => n651, Y => 
                           CARRYB_2_5_port);
   U925 : NAND2X1 port map( A => CARRYB_2_4_port, B => ab_3_4_port, Y => n652);
   U926 : NAND2X1 port map( A => ab_3_4_port, B => SUMB_2_5_port, Y => n653);
   U927 : NAND2X1 port map( A => CARRYB_2_4_port, B => SUMB_2_5_port, Y => n654
                           );
   U928 : NAND3X1 port map( A => n652, B => n653, C => n654, Y => 
                           CARRYB_3_4_port);
   U929 : NAND2X1 port map( A => SUMB_14_3_port, B => n202, Y => n655);
   U930 : NAND2X1 port map( A => SUMB_14_3_port, B => ab_15_2_port, Y => n656);
   U931 : NAND2X1 port map( A => n202, B => ab_15_2_port, Y => n657);
   U932 : NAND3X1 port map( A => n657, B => n655, C => n656, Y => 
                           CARRYB_15_2_port);
   U933 : NAND2X1 port map( A => ab_13_4_port, B => n277, Y => n658);
   U934 : NAND2X1 port map( A => SUMB_12_5_port, B => ab_13_4_port, Y => n659);
   U935 : NAND2X1 port map( A => SUMB_12_5_port, B => n277, Y => n660);
   U936 : NAND3X1 port map( A => n658, B => n659, C => n660, Y => 
                           CARRYB_13_4_port);
   U937 : NAND2X1 port map( A => ab_14_3_port, B => CARRYB_13_3_port, Y => n661
                           );
   U938 : NAND2X1 port map( A => ab_14_3_port, B => SUMB_13_4_port, Y => n662);
   U939 : NAND2X1 port map( A => CARRYB_13_3_port, B => SUMB_13_4_port, Y => 
                           n663);
   U940 : NAND3X1 port map( A => n663, B => n661, C => n662, Y => 
                           CARRYB_14_3_port);
   U941 : NAND2X1 port map( A => SUMB_5_5_port, B => n613, Y => n664);
   U942 : NAND2X1 port map( A => SUMB_5_5_port, B => ab_6_4_port, Y => n665);
   U943 : NAND2X1 port map( A => n613, B => ab_6_4_port, Y => n666);
   U944 : NAND2X1 port map( A => n41, B => n737, Y => n667);
   U945 : NAND2X1 port map( A => SUMB_1_9_port, B => n737, Y => n668);
   U946 : NAND2X1 port map( A => SUMB_1_9_port, B => n41, Y => n669);
   U947 : NAND3X1 port map( A => n667, B => n668, C => n669, Y => 
                           CARRYB_2_8_port);
   U948 : NAND2X1 port map( A => ab_3_7_port, B => CARRYB_2_7_port, Y => n670);
   U949 : NAND2X1 port map( A => SUMB_2_8_port, B => ab_3_7_port, Y => n671);
   U950 : NAND2X1 port map( A => SUMB_2_8_port, B => CARRYB_2_7_port, Y => n672
                           );
   U951 : NAND3X1 port map( A => n670, B => n671, C => n672, Y => 
                           CARRYB_3_7_port);
   U952 : NAND2X1 port map( A => SUMB_7_5_port, B => n620, Y => n673);
   U953 : NAND2X1 port map( A => SUMB_7_5_port, B => ab_8_4_port, Y => n674);
   U954 : NAND2X1 port map( A => n620, B => ab_8_4_port, Y => n675);
   U955 : NAND3X1 port map( A => n675, B => n673, C => n674, Y => 
                           CARRYB_8_4_port);
   U956 : XOR2X1 port map( A => SUMB_14_5_port, B => n676, Y => SUMB_15_4_port)
                           ;
   U957 : NAND2X1 port map( A => SUMB_14_5_port, B => n380, Y => n677);
   U958 : NAND2X1 port map( A => SUMB_14_5_port, B => ab_15_4_port, Y => n678);
   U959 : NAND2X1 port map( A => n380, B => ab_15_4_port, Y => n679);
   U960 : XOR2X1 port map( A => n680, B => SUMB_6_13_port, Y => SUMB_7_12_port)
                           ;
   U961 : NAND2X1 port map( A => ab_7_12_port, B => n713, Y => n681);
   U962 : NAND2X1 port map( A => ab_7_12_port, B => SUMB_6_13_port, Y => n682);
   U963 : NAND2X1 port map( A => n713, B => SUMB_6_13_port, Y => n683);
   U964 : NAND3X1 port map( A => n681, B => n682, C => n683, Y => 
                           CARRYB_7_12_port);
   U965 : NAND2X1 port map( A => ab_8_11_port, B => n26, Y => n684);
   U966 : NAND2X1 port map( A => ab_8_11_port, B => SUMB_7_12_port, Y => n685);
   U967 : NAND2X1 port map( A => n26, B => SUMB_7_12_port, Y => n686);
   U968 : NAND3X1 port map( A => n684, B => n685, C => n686, Y => 
                           CARRYB_8_11_port);
   U969 : XOR2X1 port map( A => ab_5_13_port, B => CARRYB_4_13_port, Y => n687)
                           ;
   U970 : XOR2X1 port map( A => n687, B => SUMB_4_14_port, Y => SUMB_5_13_port)
                           ;
   U971 : NAND2X1 port map( A => ab_5_13_port, B => CARRYB_4_13_port, Y => n688
                           );
   U972 : NAND2X1 port map( A => ab_5_13_port, B => SUMB_4_14_port, Y => n689);
   U973 : NAND2X1 port map( A => CARRYB_4_13_port, B => SUMB_4_14_port, Y => 
                           n690);
   U974 : NAND3X1 port map( A => n688, B => n689, C => n690, Y => 
                           CARRYB_5_13_port);
   U975 : NAND2X1 port map( A => ab_6_12_port, B => CARRYB_5_12_port, Y => n691
                           );
   U976 : NAND2X1 port map( A => ab_6_12_port, B => SUMB_5_13_port, Y => n692);
   U977 : NAND2X1 port map( A => CARRYB_5_12_port, B => SUMB_5_13_port, Y => 
                           n693);
   U978 : NAND3X1 port map( A => n691, B => n692, C => n693, Y => 
                           CARRYB_6_12_port);
   U979 : NAND2X1 port map( A => ab_12_7_port, B => n124, Y => n694);
   U980 : NAND2X1 port map( A => SUMB_11_8_port, B => ab_12_7_port, Y => n695);
   U981 : NAND2X1 port map( A => SUMB_11_8_port, B => n124, Y => n696);
   U982 : NAND3X1 port map( A => n694, B => n695, C => n696, Y => 
                           CARRYB_12_7_port);
   U983 : NAND2X1 port map( A => ab_13_6_port, B => n387, Y => n697);
   U984 : NAND2X1 port map( A => SUMB_12_7_port, B => ab_13_6_port, Y => n698);
   U985 : NAND2X1 port map( A => SUMB_12_7_port, B => n387, Y => n699);
   U986 : NAND3X1 port map( A => n697, B => n699, C => n698, Y => 
                           CARRYB_13_6_port);
   U987 : NAND2X1 port map( A => n245, B => ab_6_5_port, Y => n701);
   U988 : NAND2X1 port map( A => ab_6_5_port, B => SUMB_5_6_port, Y => n702);
   U989 : NAND2X1 port map( A => n245, B => SUMB_5_6_port, Y => n703);
   U990 : NAND3X1 port map( A => n701, B => n702, C => n703, Y => 
                           CARRYB_6_5_port);
   U991 : NAND2X1 port map( A => ab_7_4_port, B => n122, Y => n704);
   U992 : NAND2X1 port map( A => SUMB_6_5_port, B => ab_7_4_port, Y => n705);
   U993 : NAND2X1 port map( A => SUMB_6_5_port, B => n122, Y => n706);
   U994 : NAND3X1 port map( A => n704, B => n705, C => n706, Y => 
                           CARRYB_7_4_port);
   U995 : XOR2X1 port map( A => CARRYB_2_5_port, B => ab_3_5_port, Y => n707);
   U996 : XOR2X1 port map( A => SUMB_2_6_port, B => n707, Y => SUMB_3_5_port);
   U997 : NAND2X1 port map( A => SUMB_2_6_port, B => n533, Y => n708);
   U998 : NAND2X1 port map( A => SUMB_2_6_port, B => ab_3_5_port, Y => n709);
   U999 : NAND2X1 port map( A => n533, B => ab_3_5_port, Y => n710);
   U1000 : NAND3X1 port map( A => n709, B => n708, C => n710, Y => 
                           CARRYB_3_5_port);
   U1001 : INVX2 port map( A => CARRYB_5_12_port, Y => n711);
   U1002 : INVX2 port map( A => CARRYB_6_12_port, Y => n712);
   U1003 : BUFX4 port map( A => CARRYB_7_1_port, Y => n982);
   U1004 : NAND2X1 port map( A => ab_9_6_port, B => n442, Y => n714);
   U1005 : NAND2X1 port map( A => SUMB_8_7_port, B => ab_9_6_port, Y => n715);
   U1006 : NAND2X1 port map( A => SUMB_8_7_port, B => n442, Y => n716);
   U1007 : NAND3X1 port map( A => n714, B => n715, C => n716, Y => 
                           CARRYB_9_6_port);
   U1008 : NAND2X1 port map( A => n179, B => ab_10_5_port, Y => n717);
   U1009 : NAND2X1 port map( A => SUMB_9_6_port, B => n179, Y => n718);
   U1010 : NAND2X1 port map( A => SUMB_9_6_port, B => ab_10_5_port, Y => n719);
   U1011 : NAND3X1 port map( A => n717, B => n718, C => n719, Y => 
                           CARRYB_10_5_port);
   U1012 : XOR2X1 port map( A => A(15), B => B(15), Y => n720);
   U1013 : XOR2X1 port map( A => n315, B => n720, Y => A1_13_port);
   U1014 : NAND2X1 port map( A => SUMB_15_0_port, B => A(15), Y => n721);
   U1015 : NAND2X1 port map( A => SUMB_15_0_port, B => B(15), Y => n722);
   U1016 : NAND2X1 port map( A => A(15), B => B(15), Y => n723);
   U1017 : NAND3X1 port map( A => n723, B => n721, C => n722, Y => A2_14_port);
   U1018 : XNOR2X1 port map( A => n724, B => SUMB_9_2_port, Y => SUMB_10_1_port
                           );
   U1019 : XNOR2X1 port map( A => n433, B => ab_10_1_port, Y => n724);
   U1020 : XOR2X1 port map( A => ab_5_10_port, B => CARRYB_4_10_port, Y => n725
                           );
   U1021 : NAND2X1 port map( A => ab_5_10_port, B => CARRYB_4_10_port, Y => 
                           n727);
   U1022 : NAND2X1 port map( A => ab_5_10_port, B => SUMB_4_11_port, Y => n728)
                           ;
   U1023 : NAND2X1 port map( A => CARRYB_4_10_port, B => SUMB_4_11_port, Y => 
                           n729);
   U1024 : NAND3X1 port map( A => n727, B => n728, C => n729, Y => 
                           CARRYB_5_10_port);
   U1025 : NAND2X1 port map( A => ab_6_9_port, B => CARRYB_5_9_port, Y => n730)
                           ;
   U1026 : NAND2X1 port map( A => ab_6_9_port, B => SUMB_5_10_port, Y => n731);
   U1027 : NAND2X1 port map( A => CARRYB_5_9_port, B => SUMB_5_10_port, Y => 
                           n732);
   U1028 : NAND3X1 port map( A => n730, B => n731, C => n732, Y => 
                           CARRYB_6_9_port);
   U1029 : NAND2X1 port map( A => SUMB_3_12_port, B => n348, Y => n733);
   U1030 : NAND2X1 port map( A => SUMB_3_12_port, B => ab_4_11_port, Y => n734)
                           ;
   U1031 : NAND2X1 port map( A => n348, B => ab_4_11_port, Y => n735);
   U1032 : NAND3X1 port map( A => n735, B => n734, C => n733, Y => 
                           CARRYB_4_11_port);
   U1033 : BUFX2 port map( A => CARRYB_4_8_port, Y => n981);
   U1034 : XNOR2X1 port map( A => n960, B => ab_7_2_port, Y => n930);
   U1035 : INVX2 port map( A => B(1), Y => n992);
   U1036 : NAND2X1 port map( A => ab_3_13_port, B => n60, Y => n738);
   U1037 : NAND2X1 port map( A => ab_3_13_port, B => SUMB_2_14_port, Y => n739)
                           ;
   U1038 : NAND2X1 port map( A => n60, B => SUMB_2_14_port, Y => n740);
   U1039 : NAND3X1 port map( A => n738, B => n739, C => n740, Y => 
                           CARRYB_3_13_port);
   U1040 : NAND2X1 port map( A => ab_4_12_port, B => n594, Y => n741);
   U1041 : NAND2X1 port map( A => SUMB_3_13_port, B => ab_4_12_port, Y => n742)
                           ;
   U1042 : NAND2X1 port map( A => n594, B => SUMB_3_13_port, Y => n743);
   U1043 : NAND3X1 port map( A => n741, B => n742, C => n743, Y => 
                           CARRYB_4_12_port);
   U1044 : NAND2X1 port map( A => ab_9_8_port, B => n388, Y => n744);
   U1045 : NAND2X1 port map( A => ab_9_8_port, B => SUMB_8_9_port, Y => n745);
   U1046 : NAND2X1 port map( A => n388, B => SUMB_8_9_port, Y => n746);
   U1047 : NAND3X1 port map( A => n744, B => n745, C => n746, Y => 
                           CARRYB_9_8_port);
   U1048 : NAND2X1 port map( A => ab_10_7_port, B => n539, Y => n747);
   U1049 : NAND2X1 port map( A => ab_10_7_port, B => SUMB_9_8_port, Y => n748);
   U1050 : NAND2X1 port map( A => n539, B => SUMB_9_8_port, Y => n749);
   U1051 : NAND3X1 port map( A => n747, B => n748, C => n749, Y => 
                           CARRYB_10_7_port);
   U1052 : XNOR2X1 port map( A => n750, B => SUMB_6_11_port, Y => 
                           SUMB_7_10_port);
   U1053 : XOR2X1 port map( A => SUMB_7_3_port, B => ab_8_2_port, Y => n751);
   U1054 : XOR2X1 port map( A => n751, B => n92, Y => SUMB_8_2_port);
   U1055 : NAND2X1 port map( A => SUMB_11_2_port, B => CARRYB_11_1_port, Y => 
                           n752);
   U1056 : NAND2X1 port map( A => CARRYB_11_1_port, B => ab_12_1_port, Y => 
                           n753);
   U1057 : NAND2X1 port map( A => SUMB_11_2_port, B => ab_12_1_port, Y => n754)
                           ;
   U1058 : NAND3X1 port map( A => n753, B => n754, C => n752, Y => 
                           CARRYB_12_1_port);
   U1059 : NAND2X1 port map( A => SUMB_5_8_port, B => CARRYB_5_7_port, Y => 
                           n756);
   U1060 : NAND2X1 port map( A => CARRYB_5_7_port, B => ab_6_7_port, Y => n757)
                           ;
   U1061 : NAND2X1 port map( A => SUMB_5_8_port, B => ab_6_7_port, Y => n758);
   U1062 : NAND3X1 port map( A => n758, B => n756, C => n757, Y => 
                           CARRYB_6_7_port);
   U1063 : XOR2X1 port map( A => n260, B => ab_5_4_port, Y => n759);
   U1064 : XOR2X1 port map( A => n121, B => n759, Y => SUMB_5_4_port);
   U1065 : NAND2X1 port map( A => SUMB_4_5_port, B => n260, Y => n760);
   U1066 : NAND2X1 port map( A => SUMB_4_5_port, B => ab_5_4_port, Y => n761);
   U1067 : NAND2X1 port map( A => n260, B => ab_5_4_port, Y => n762);
   U1068 : NAND3X1 port map( A => n761, B => n762, C => n760, Y => 
                           CARRYB_5_4_port);
   U1069 : NAND2X1 port map( A => ab_10_4_port, B => n38, Y => n764);
   U1070 : NAND2X1 port map( A => SUMB_9_5_port, B => ab_10_4_port, Y => n765);
   U1071 : NAND2X1 port map( A => SUMB_9_5_port, B => n38, Y => n766);
   U1072 : NAND3X1 port map( A => n764, B => n765, C => n766, Y => 
                           CARRYB_10_4_port);
   U1073 : NAND2X1 port map( A => ab_11_3_port, B => n484, Y => n767);
   U1074 : NAND2X1 port map( A => ab_11_3_port, B => SUMB_10_4_port, Y => n768)
                           ;
   U1075 : NAND2X1 port map( A => SUMB_10_4_port, B => n484, Y => n769);
   U1076 : NAND3X1 port map( A => n767, B => n768, C => n769, Y => 
                           CARRYB_11_3_port);
   U1077 : XOR2X1 port map( A => n313, B => ab_7_11_port, Y => n770);
   U1078 : XOR2X1 port map( A => n770, B => n117, Y => SUMB_7_11_port);
   U1079 : XOR2X1 port map( A => CARRYB_7_10_port, B => ab_8_10_port, Y => n771
                           );
   U1080 : XOR2X1 port map( A => n771, B => SUMB_7_11_port, Y => SUMB_8_10_port
                           );
   U1081 : NAND2X1 port map( A => ab_7_11_port, B => CARRYB_6_11_port, Y => 
                           n772);
   U1082 : NAND2X1 port map( A => ab_7_11_port, B => SUMB_6_12_port, Y => n773)
                           ;
   U1083 : NAND2X1 port map( A => CARRYB_6_11_port, B => SUMB_6_12_port, Y => 
                           n774);
   U1084 : NAND3X1 port map( A => n772, B => n773, C => n774, Y => 
                           CARRYB_7_11_port);
   U1085 : NAND2X1 port map( A => ab_8_10_port, B => CARRYB_7_10_port, Y => 
                           n775);
   U1086 : NAND2X1 port map( A => ab_8_10_port, B => SUMB_7_11_port, Y => n776)
                           ;
   U1087 : NAND2X1 port map( A => CARRYB_7_10_port, B => SUMB_7_11_port, Y => 
                           n777);
   U1088 : NAND3X1 port map( A => n775, B => n776, C => n777, Y => 
                           CARRYB_8_10_port);
   U1089 : NAND2X1 port map( A => ab_13_5_port, B => n540, Y => n778);
   U1090 : NAND2X1 port map( A => SUMB_12_6_port, B => ab_13_5_port, Y => n779)
                           ;
   U1091 : NAND2X1 port map( A => SUMB_12_6_port, B => n540, Y => n780);
   U1092 : NAND3X1 port map( A => n778, B => n779, C => n780, Y => 
                           CARRYB_13_5_port);
   U1093 : NAND2X1 port map( A => ab_14_4_port, B => n330, Y => n781);
   U1094 : NAND2X1 port map( A => SUMB_13_5_port, B => ab_14_4_port, Y => n782)
                           ;
   U1095 : NAND2X1 port map( A => SUMB_13_5_port, B => n330, Y => n783);
   U1096 : NAND3X1 port map( A => n781, B => n783, C => n782, Y => 
                           CARRYB_14_4_port);
   U1097 : NAND2X1 port map( A => ab_8_8_port, B => n278, Y => n784);
   U1098 : NAND2X1 port map( A => SUMB_7_9_port, B => ab_8_8_port, Y => n785);
   U1099 : NAND2X1 port map( A => n278, B => SUMB_7_9_port, Y => n786);
   U1100 : NAND3X1 port map( A => n784, B => n785, C => n786, Y => 
                           CARRYB_8_8_port);
   U1101 : NAND2X1 port map( A => ab_9_7_port, B => n381, Y => n787);
   U1102 : NAND2X1 port map( A => SUMB_8_8_port, B => ab_9_7_port, Y => n788);
   U1103 : NAND2X1 port map( A => SUMB_8_8_port, B => n381, Y => n789);
   U1104 : NAND3X1 port map( A => n787, B => n788, C => n789, Y => 
                           CARRYB_9_7_port);
   U1105 : XOR2X1 port map( A => ab_6_10_port, B => CARRYB_5_10_port, Y => n790
                           );
   U1106 : XOR2X1 port map( A => n790, B => n95, Y => SUMB_6_10_port);
   U1107 : XOR2X1 port map( A => ab_7_9_port, B => CARRYB_6_9_port, Y => n791);
   U1108 : NAND2X1 port map( A => ab_6_10_port, B => CARRYB_5_10_port, Y => 
                           n792);
   U1109 : NAND2X1 port map( A => SUMB_5_11_port, B => ab_6_10_port, Y => n793)
                           ;
   U1110 : NAND2X1 port map( A => SUMB_5_11_port, B => CARRYB_5_10_port, Y => 
                           n794);
   U1111 : NAND3X1 port map( A => n792, B => n793, C => n794, Y => 
                           CARRYB_6_10_port);
   U1112 : NAND2X1 port map( A => ab_7_9_port, B => n56, Y => n795);
   U1113 : NAND2X1 port map( A => ab_7_9_port, B => SUMB_6_10_port, Y => n796);
   U1114 : NAND2X1 port map( A => n56, B => SUMB_6_10_port, Y => n797);
   U1115 : NAND3X1 port map( A => n795, B => n796, C => n797, Y => 
                           CARRYB_7_9_port);
   U1116 : NAND2X1 port map( A => n811, B => n79, Y => n979);
   U1117 : NAND2X1 port map( A => SUMB_10_2_port, B => n84, Y => n798);
   U1118 : NAND2X1 port map( A => SUMB_10_2_port, B => ab_11_1_port, Y => n799)
                           ;
   U1119 : NAND2X1 port map( A => n84, B => ab_11_1_port, Y => n800);
   U1120 : NAND3X1 port map( A => n799, B => n800, C => n798, Y => 
                           CARRYB_11_1_port);
   U1121 : NAND2X1 port map( A => SUMB_6_4_port, B => CARRYB_6_3_port, Y => 
                           n801);
   U1122 : NAND2X1 port map( A => SUMB_6_4_port, B => ab_7_3_port, Y => n802);
   U1123 : NAND2X1 port map( A => CARRYB_6_3_port, B => ab_7_3_port, Y => n803)
                           ;
   U1124 : NAND3X1 port map( A => n803, B => n802, C => n801, Y => 
                           CARRYB_7_3_port);
   U1125 : NAND2X1 port map( A => ab_6_11_port, B => CARRYB_5_11_port, Y => 
                           n804);
   U1126 : NAND2X1 port map( A => ab_6_11_port, B => SUMB_5_12_port, Y => n805)
                           ;
   U1127 : NAND2X1 port map( A => CARRYB_5_11_port, B => SUMB_5_12_port, Y => 
                           n806);
   U1128 : NAND3X1 port map( A => n804, B => n805, C => n806, Y => 
                           CARRYB_6_11_port);
   U1129 : NAND2X1 port map( A => ab_7_10_port, B => n557, Y => n807);
   U1130 : NAND2X1 port map( A => ab_7_10_port, B => SUMB_6_11_port, Y => n808)
                           ;
   U1131 : NAND2X1 port map( A => SUMB_6_11_port, B => n557, Y => n809);
   U1132 : NAND3X1 port map( A => n807, B => n808, C => n809, Y => 
                           CARRYB_7_10_port);
   U1133 : NAND2X1 port map( A => n173, B => SUMB_7_4_port, Y => n810);
   U1134 : NAND2X1 port map( A => SUMB_7_4_port, B => ab_8_3_port, Y => n811);
   U1135 : NAND2X1 port map( A => n173, B => ab_8_3_port, Y => n812);
   U1136 : NAND3X1 port map( A => n811, B => n812, C => n810, Y => 
                           CARRYB_8_3_port);
   U1137 : INVX2 port map( A => A(1), Y => n986);
   U1138 : NAND2X1 port map( A => SUMB_3_10_port, B => n978, Y => n813);
   U1139 : NAND2X1 port map( A => n978, B => ab_4_9_port, Y => n814);
   U1140 : NAND2X1 port map( A => SUMB_3_10_port, B => ab_4_9_port, Y => n815);
   U1141 : NAND3X1 port map( A => n814, B => n813, C => n815, Y => 
                           CARRYB_4_9_port);
   U1142 : NAND2X1 port map( A => SUMB_1_11_port, B => n77, Y => n816);
   U1143 : NAND2X1 port map( A => n77, B => ab_2_10_port, Y => n817);
   U1144 : NAND2X1 port map( A => SUMB_1_11_port, B => ab_2_10_port, Y => n818)
                           ;
   U1145 : NAND3X1 port map( A => n817, B => n816, C => n818, Y => 
                           CARRYB_2_10_port);
   U1146 : NAND2X1 port map( A => ab_4_6_port, B => n246, Y => n819);
   U1147 : NAND2X1 port map( A => SUMB_3_7_port, B => ab_4_6_port, Y => n820);
   U1148 : NAND2X1 port map( A => n246, B => SUMB_3_7_port, Y => n821);
   U1149 : NAND3X1 port map( A => n819, B => n820, C => n821, Y => 
                           CARRYB_4_6_port);
   U1150 : NAND2X1 port map( A => ab_5_5_port, B => n523, Y => n822);
   U1151 : NAND2X1 port map( A => SUMB_4_6_port, B => ab_5_5_port, Y => n823);
   U1152 : NAND2X1 port map( A => SUMB_4_6_port, B => n523, Y => n824);
   U1153 : NAND3X1 port map( A => n824, B => n822, C => n823, Y => 
                           CARRYB_5_5_port);
   U1154 : NAND2X1 port map( A => n435, B => n61, Y => n825);
   U1155 : NAND2X1 port map( A => SUMB_1_8_port, B => n435, Y => n826);
   U1156 : NAND2X1 port map( A => n61, B => SUMB_1_8_port, Y => n827);
   U1157 : NAND3X1 port map( A => n825, B => n826, C => n827, Y => 
                           CARRYB_2_7_port);
   U1158 : NAND2X1 port map( A => n848, B => ab_3_6_port, Y => n828);
   U1159 : NAND2X1 port map( A => SUMB_2_7_port, B => ab_3_6_port, Y => n829);
   U1160 : NAND2X1 port map( A => n848, B => SUMB_2_7_port, Y => n830);
   U1161 : NAND3X1 port map( A => n829, B => n828, C => n830, Y => 
                           CARRYB_3_6_port);
   U1162 : NAND2X1 port map( A => SUMB_6_6_port, B => CARRYB_6_5_port, Y => 
                           n831);
   U1163 : NAND2X1 port map( A => CARRYB_6_5_port, B => ab_7_5_port, Y => n832)
                           ;
   U1164 : NAND2X1 port map( A => SUMB_6_6_port, B => ab_7_5_port, Y => n833);
   U1165 : NAND3X1 port map( A => n832, B => n831, C => n833, Y => 
                           CARRYB_7_5_port);
   U1166 : NAND2X1 port map( A => ab_8_5_port, B => n303, Y => n834);
   U1167 : NAND2X1 port map( A => SUMB_7_6_port, B => ab_8_5_port, Y => n835);
   U1168 : NAND2X1 port map( A => SUMB_7_6_port, B => n303, Y => n836);
   U1169 : NAND3X1 port map( A => n834, B => n835, C => n836, Y => 
                           CARRYB_8_5_port);
   U1170 : NAND2X1 port map( A => n98, B => ab_9_4_port, Y => n837);
   U1171 : NAND2X1 port map( A => SUMB_8_5_port, B => n98, Y => n838);
   U1172 : NAND2X1 port map( A => SUMB_8_5_port, B => ab_9_4_port, Y => n839);
   U1173 : NAND3X1 port map( A => n837, B => n839, C => n838, Y => 
                           CARRYB_9_4_port);
   U1174 : NAND2X1 port map( A => ab_3_8_port, B => n126, Y => n840);
   U1175 : NAND2X1 port map( A => SUMB_2_9_port, B => ab_3_8_port, Y => n841);
   U1176 : NAND2X1 port map( A => SUMB_2_9_port, B => n126, Y => n842);
   U1177 : NAND3X1 port map( A => n840, B => n841, C => n842, Y => 
                           CARRYB_3_8_port);
   U1178 : NAND2X1 port map( A => ab_4_7_port, B => n494, Y => n843);
   U1179 : NAND2X1 port map( A => SUMB_3_8_port, B => ab_4_7_port, Y => n844);
   U1180 : NAND2X1 port map( A => SUMB_3_8_port, B => n494, Y => n845);
   U1181 : NAND3X1 port map( A => n843, B => n844, C => n845, Y => 
                           CARRYB_4_7_port);
   U1182 : INVX2 port map( A => CARRYB_2_6_port, Y => n847);
   U1183 : XOR2X1 port map( A => n164, B => ab_9_0_port, Y => n849);
   U1184 : XOR2X1 port map( A => CARRYB_8_0_port, B => n849, Y => A1_7_port);
   U1185 : NAND2X1 port map( A => SUMB_8_1_port, B => CARRYB_8_0_port, Y => 
                           n850);
   U1186 : NAND2X1 port map( A => CARRYB_8_0_port, B => ab_9_0_port, Y => n851)
                           ;
   U1187 : NAND2X1 port map( A => SUMB_8_1_port, B => ab_9_0_port, Y => n852);
   U1188 : NAND3X1 port map( A => n851, B => n850, C => n852, Y => 
                           CARRYB_9_0_port);
   U1189 : XOR2X1 port map( A => n344, B => ab_10_0_port, Y => n853);
   U1190 : XOR2X1 port map( A => n89, B => n853, Y => A1_8_port);
   U1191 : NAND2X1 port map( A => SUMB_9_1_port, B => CARRYB_9_0_port, Y => 
                           n854);
   U1192 : NAND2X1 port map( A => SUMB_9_1_port, B => ab_10_0_port, Y => n855);
   U1193 : NAND2X1 port map( A => CARRYB_9_0_port, B => ab_10_0_port, Y => n856
                           );
   U1194 : NAND3X1 port map( A => n855, B => n856, C => n854, Y => 
                           CARRYB_10_0_port);
   U1195 : XOR2X1 port map( A => n857, B => SUMB_4_2_port, Y => SUMB_5_1_port);
   U1196 : NAND2X1 port map( A => SUMB_4_2_port, B => CARRYB_4_1_port, Y => 
                           n858);
   U1197 : NAND2X1 port map( A => SUMB_4_2_port, B => ab_5_1_port, Y => n859);
   U1198 : NAND2X1 port map( A => CARRYB_4_1_port, B => ab_5_1_port, Y => n860)
                           ;
   U1199 : NAND3X1 port map( A => n859, B => n858, C => n860, Y => 
                           CARRYB_5_1_port);
   U1200 : XOR2X1 port map( A => ab_7_0_port, B => n989, Y => n861);
   U1201 : XOR2X1 port map( A => n861, B => SUMB_6_1_port, Y => A1_5_port);
   U1202 : NAND2X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, Y => n862)
                           ;
   U1203 : NAND2X1 port map( A => ab_6_1_port, B => SUMB_5_2_port, Y => n863);
   U1204 : NAND2X1 port map( A => CARRYB_5_1_port, B => SUMB_5_2_port, Y => 
                           n864);
   U1205 : NAND3X1 port map( A => n862, B => n863, C => n864, Y => 
                           CARRYB_6_1_port);
   U1206 : NAND2X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, Y => n865)
                           ;
   U1207 : NAND2X1 port map( A => ab_7_0_port, B => SUMB_6_1_port, Y => n866);
   U1208 : NAND2X1 port map( A => CARRYB_6_0_port, B => SUMB_6_1_port, Y => 
                           n867);
   U1209 : NAND3X1 port map( A => n865, B => n866, C => n867, Y => 
                           CARRYB_7_0_port);
   U1210 : XOR2X1 port map( A => CARRYB_3_2_port, B => ab_4_2_port, Y => n868);
   U1211 : XOR2X1 port map( A => n627, B => n868, Y => SUMB_4_2_port);
   U1212 : NAND2X1 port map( A => SUMB_3_3_port, B => n190, Y => n869);
   U1213 : NAND2X1 port map( A => SUMB_3_3_port, B => ab_4_2_port, Y => n870);
   U1214 : NAND2X1 port map( A => n190, B => ab_4_2_port, Y => n871);
   U1215 : NAND3X1 port map( A => n870, B => n869, C => n871, Y => 
                           CARRYB_4_2_port);
   U1216 : NAND2X1 port map( A => CARRYB_1_12_port, B => ab_2_12_port, Y => 
                           n872);
   U1217 : NAND2X1 port map( A => CARRYB_1_12_port, B => SUMB_1_13_port, Y => 
                           n873);
   U1218 : NAND2X1 port map( A => ab_2_12_port, B => SUMB_1_13_port, Y => n874)
                           ;
   U1219 : NAND3X1 port map( A => n872, B => n873, C => n874, Y => 
                           CARRYB_2_12_port);
   U1220 : NAND2X1 port map( A => ab_3_11_port, B => n385, Y => n875);
   U1221 : NAND2X1 port map( A => SUMB_2_12_port, B => ab_3_11_port, Y => n876)
                           ;
   U1222 : NAND2X1 port map( A => SUMB_2_12_port, B => n385, Y => n877);
   U1223 : NAND3X1 port map( A => n875, B => n876, C => n877, Y => 
                           CARRYB_3_11_port);
   U1224 : NAND2X1 port map( A => ab_7_8_port, B => n299, Y => n878);
   U1225 : NAND2X1 port map( A => SUMB_6_9_port, B => ab_7_8_port, Y => n879);
   U1226 : NAND2X1 port map( A => SUMB_6_9_port, B => n299, Y => n880);
   U1227 : NAND3X1 port map( A => n878, B => n879, C => n880, Y => 
                           CARRYB_7_8_port);
   U1228 : NAND2X1 port map( A => ab_8_7_port, B => n329, Y => n881);
   U1229 : NAND2X1 port map( A => SUMB_7_8_port, B => ab_8_7_port, Y => n882);
   U1230 : NAND2X1 port map( A => SUMB_7_8_port, B => n329, Y => n883);
   U1231 : NAND3X1 port map( A => n881, B => n882, C => n883, Y => 
                           CARRYB_8_7_port);
   U1232 : NAND2X1 port map( A => ab_9_2_port, B => CARRYB_8_2_port, Y => n884)
                           ;
   U1233 : NAND2X1 port map( A => SUMB_8_3_port, B => ab_9_2_port, Y => n885);
   U1234 : NAND2X1 port map( A => CARRYB_8_2_port, B => SUMB_8_3_port, Y => 
                           n886);
   U1235 : NAND3X1 port map( A => n885, B => n884, C => n886, Y => 
                           CARRYB_9_2_port);
   U1236 : NAND2X1 port map( A => CARRYB_9_1_port, B => ab_10_1_port, Y => n887
                           );
   U1237 : NAND2X1 port map( A => SUMB_9_2_port, B => CARRYB_9_1_port, Y => 
                           n888);
   U1238 : NAND2X1 port map( A => ab_10_1_port, B => SUMB_9_2_port, Y => n889);
   U1239 : NAND3X1 port map( A => n887, B => n888, C => n889, Y => 
                           CARRYB_10_1_port);
   U1240 : NAND2X1 port map( A => SUMB_4_10_port, B => n378, Y => n890);
   U1241 : NAND2X1 port map( A => SUMB_4_10_port, B => ab_5_9_port, Y => n891);
   U1242 : NAND2X1 port map( A => n378, B => ab_5_9_port, Y => n892);
   U1243 : NAND3X1 port map( A => n891, B => n892, C => n890, Y => 
                           CARRYB_5_9_port);
   U1244 : NAND2X1 port map( A => ab_6_8_port, B => n490, Y => n893);
   U1245 : NAND2X1 port map( A => SUMB_5_9_port, B => ab_6_8_port, Y => n894);
   U1246 : NAND2X1 port map( A => SUMB_5_9_port, B => n490, Y => n895);
   U1247 : NAND3X1 port map( A => n893, B => n894, C => n895, Y => 
                           CARRYB_6_8_port);
   U1248 : NAND2X1 port map( A => ab_7_7_port, B => n488, Y => n896);
   U1249 : NAND2X1 port map( A => SUMB_6_8_port, B => ab_7_7_port, Y => n897);
   U1250 : NAND2X1 port map( A => SUMB_6_8_port, B => n488, Y => n898);
   U1251 : NAND3X1 port map( A => n896, B => n897, C => n898, Y => 
                           CARRYB_7_7_port);
   U1252 : NAND2X1 port map( A => n222, B => ab_2_11_port, Y => n899);
   U1253 : NAND2X1 port map( A => n222, B => SUMB_1_12_port, Y => n900);
   U1254 : NAND2X1 port map( A => ab_2_11_port, B => SUMB_1_12_port, Y => n901)
                           ;
   U1255 : NAND3X1 port map( A => n899, B => n900, C => n901, Y => 
                           CARRYB_2_11_port);
   U1256 : NAND2X1 port map( A => ab_3_10_port, B => n910, Y => n902);
   U1257 : NAND2X1 port map( A => n223, B => ab_3_10_port, Y => n903);
   U1258 : NAND2X1 port map( A => n223, B => n910, Y => n904);
   U1259 : NAND3X1 port map( A => n902, B => n904, C => n903, Y => 
                           CARRYB_3_10_port);
   U1260 : INVX2 port map( A => CARRYB_3_0_port, Y => n905);
   U1261 : INVX4 port map( A => n905, Y => n906);
   U1262 : INVX2 port map( A => CARRYB_4_0_port, Y => n907);
   U1263 : INVX4 port map( A => n907, Y => n908);
   U1264 : NAND2X1 port map( A => SUMB_8_4_port, B => n979, Y => n911);
   U1265 : NAND2X1 port map( A => SUMB_8_4_port, B => ab_9_3_port, Y => n912);
   U1266 : NAND2X1 port map( A => n979, B => ab_9_3_port, Y => n913);
   U1267 : NAND3X1 port map( A => n913, B => n912, C => n911, Y => 
                           CARRYB_9_3_port);
   U1268 : NAND2X1 port map( A => n491, B => ab_10_3_port, Y => n914);
   U1269 : NAND2X1 port map( A => SUMB_9_4_port, B => ab_10_3_port, Y => n915);
   U1270 : NAND2X1 port map( A => SUMB_9_4_port, B => n491, Y => n916);
   U1271 : NAND3X1 port map( A => n914, B => n915, C => n916, Y => 
                           CARRYB_10_3_port);
   U1272 : NAND2X1 port map( A => n85, B => ab_11_2_port, Y => n917);
   U1273 : NAND2X1 port map( A => SUMB_10_3_port, B => ab_11_2_port, Y => n918)
                           ;
   U1274 : NAND2X1 port map( A => SUMB_10_3_port, B => n85, Y => n919);
   U1275 : NAND3X1 port map( A => n917, B => n918, C => n919, Y => 
                           CARRYB_11_2_port);
   U1276 : NAND2X1 port map( A => SUMB_2_10_port, B => n977, Y => n920);
   U1277 : NAND2X1 port map( A => SUMB_2_10_port, B => ab_3_9_port, Y => n921);
   U1278 : NAND2X1 port map( A => n977, B => ab_3_9_port, Y => n922);
   U1279 : NAND3X1 port map( A => n922, B => n920, C => n921, Y => 
                           CARRYB_3_9_port);
   U1280 : XOR2X1 port map( A => n923, B => SUMB_5_7_port, Y => SUMB_6_6_port);
   U1281 : NAND2X1 port map( A => ab_5_7_port, B => n270, Y => n924);
   U1282 : NAND2X1 port map( A => n247, B => ab_5_7_port, Y => n925);
   U1283 : NAND2X1 port map( A => n247, B => n270, Y => n926);
   U1284 : NAND3X1 port map( A => n924, B => n925, C => n926, Y => 
                           CARRYB_5_7_port);
   U1285 : NAND2X1 port map( A => n193, B => ab_6_6_port, Y => n927);
   U1286 : NAND2X1 port map( A => SUMB_5_7_port, B => ab_6_6_port, Y => n928);
   U1287 : NAND2X1 port map( A => SUMB_5_7_port, B => n230, Y => n929);
   U1288 : NAND3X1 port map( A => n927, B => n929, C => n928, Y => 
                           CARRYB_6_6_port);
   U1289 : XOR2X1 port map( A => n930, B => n531, Y => SUMB_7_2_port);
   U1290 : XOR2X1 port map( A => ab_8_1_port, B => n982, Y => n931);
   U1291 : NAND2X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, Y => n932)
                           ;
   U1292 : NAND2X1 port map( A => ab_7_2_port, B => SUMB_6_3_port, Y => n933);
   U1293 : NAND2X1 port map( A => CARRYB_6_2_port, B => SUMB_6_3_port, Y => 
                           n934);
   U1294 : NAND3X1 port map( A => n932, B => n933, C => n934, Y => 
                           CARRYB_7_2_port);
   U1295 : NAND2X1 port map( A => ab_8_1_port, B => n982, Y => n935);
   U1296 : NAND2X1 port map( A => ab_8_1_port, B => SUMB_7_2_port, Y => n936);
   U1297 : NAND2X1 port map( A => n982, B => SUMB_7_2_port, Y => n937);
   U1298 : NAND3X1 port map( A => n936, B => n935, C => n937, Y => 
                           CARRYB_8_1_port);
   U1299 : NAND2X1 port map( A => CARRYB_2_3_port, B => n951, Y => n940);
   U1300 : NAND2X1 port map( A => n938, B => n939, Y => n941);
   U1301 : NAND2X1 port map( A => n940, B => n941, Y => SUMB_3_3_port);
   U1302 : INVX1 port map( A => CARRYB_2_3_port, Y => n938);
   U1303 : NAND2X1 port map( A => SUMB_6_7_port, B => n614, Y => n942);
   U1304 : NAND2X1 port map( A => SUMB_6_7_port, B => ab_7_6_port, Y => n943);
   U1305 : NAND2X1 port map( A => n614, B => ab_7_6_port, Y => n944);
   U1306 : NAND3X1 port map( A => n944, B => n943, C => n942, Y => 
                           CARRYB_7_6_port);
   U1307 : XOR2X1 port map( A => CARRYB_4_8_port, B => ab_5_8_port, Y => n945);
   U1308 : XOR2X1 port map( A => SUMB_4_9_port, B => n945, Y => SUMB_5_8_port);
   U1309 : NAND2X1 port map( A => SUMB_4_9_port, B => n981, Y => n946);
   U1310 : NAND2X1 port map( A => SUMB_4_9_port, B => ab_5_8_port, Y => n947);
   U1311 : NAND2X1 port map( A => n981, B => ab_5_8_port, Y => n948);
   U1312 : NAND3X1 port map( A => n948, B => n947, C => n946, Y => 
                           CARRYB_5_8_port);
   U1313 : AND2X2 port map( A => n524, B => ab_1_5_port, Y => n950);
   U1314 : INVX4 port map( A => A(2), Y => n1022);
   U1315 : XNOR2X1 port map( A => SUMB_2_4_port, B => ab_3_3_port, Y => n951);
   U1316 : INVX2 port map( A => CARRYB_4_1_port, Y => n952);
   U1317 : XOR2X1 port map( A => CARRYB_2_2_port, B => ab_3_2_port, Y => n953);
   U1318 : XOR2X1 port map( A => SUMB_2_3_port, B => n953, Y => SUMB_3_2_port);
   U1319 : NAND2X1 port map( A => SUMB_2_3_port, B => CARRYB_2_2_port, Y => 
                           n954);
   U1320 : NAND2X1 port map( A => SUMB_2_3_port, B => ab_3_2_port, Y => n955);
   U1321 : NAND2X1 port map( A => CARRYB_2_2_port, B => ab_3_2_port, Y => n956)
                           ;
   U1322 : NAND3X1 port map( A => n955, B => n954, C => n956, Y => 
                           CARRYB_3_2_port);
   U1323 : NAND2X1 port map( A => SUMB_7_3_port, B => CARRYB_7_2_port, Y => 
                           n957);
   U1324 : NAND2X1 port map( A => CARRYB_7_2_port, B => ab_8_2_port, Y => n958)
                           ;
   U1325 : NAND2X1 port map( A => SUMB_7_3_port, B => ab_8_2_port, Y => n959);
   U1326 : NAND3X1 port map( A => n959, B => n957, C => n958, Y => 
                           CARRYB_8_2_port);
   U1327 : NAND2X1 port map( A => CARRYB_2_3_port, B => SUMB_2_4_port, Y => 
                           n961);
   U1328 : NAND2X1 port map( A => CARRYB_2_3_port, B => ab_3_3_port, Y => n962)
                           ;
   U1329 : NAND2X1 port map( A => ab_3_3_port, B => SUMB_2_4_port, Y => n963);
   U1330 : NAND3X1 port map( A => n962, B => n963, C => n961, Y => 
                           CARRYB_3_3_port);
   U1331 : AND2X2 port map( A => CARRYB_15_0_port, B => SUMB_15_1_port, Y => 
                           n972);
   U1332 : AND2X2 port map( A => n1025, B => n1009, Y => ab_3_9_port);
   U1333 : NOR2X1 port map( A => n1021, B => n994, Y => n964);
   U1334 : INVX1 port map( A => CARRYB_6_0_port, Y => n988);
   U1335 : AND2X2 port map( A => ab_0_5_port, B => n525, Y => n965);
   U1336 : AND2X2 port map( A => n228, B => CARRYB_15_4_port, Y => n968);
   U1337 : AND2X2 port map( A => ab_0_2_port, B => ab_1_1_port, Y => n969);
   U1338 : AND2X2 port map( A => ab_1_3_port, B => ab_0_4_port, Y => n970);
   U1339 : AND2X2 port map( A => SUMB_15_6_port, B => CARRYB_15_5_port, Y => 
                           n973);
   U1340 : INVX4 port map( A => n992, Y => n993);
   U1341 : INVX2 port map( A => n988, Y => n989);
   U1342 : INVX2 port map( A => B(0), Y => n990);
   U1343 : INVX2 port map( A => A(13), Y => n1052);
   U1344 : INVX2 port map( A => A(15), Y => n1050);
   U1345 : INVX2 port map( A => A(14), Y => n1051);
   U1346 : INVX2 port map( A => A(4), Y => n1026);
   U1347 : INVX2 port map( A => A(6), Y => n1030);
   U1348 : INVX2 port map( A => A(5), Y => n1028);
   U1349 : INVX2 port map( A => A(8), Y => n1034);
   U1350 : INVX2 port map( A => A(7), Y => n1032);
   U1351 : INVX2 port map( A => A(9), Y => n1036);
   U1352 : XOR2X1 port map( A => CARRYB_15_0_port, B => SUMB_15_1_port, Y => 
                           A1_14_port);
   U1353 : XOR2X1 port map( A => CARRYB_15_1_port, B => SUMB_15_2_port, Y => 
                           A1_15_port);
   U1354 : XOR2X1 port map( A => SUMB_15_3_port, B => CARRYB_15_2_port, Y => 
                           A1_16_port);
   U1355 : XOR2X1 port map( A => SUMB_15_4_port, B => CARRYB_15_3_port, Y => 
                           A1_17_port);
   U1356 : XOR2X1 port map( A => SUMB_15_7_port, B => CARRYB_15_6_port, Y => 
                           A1_20_port);
   U1357 : XOR2X1 port map( A => SUMB_15_8_port, B => CARRYB_15_7_port, Y => 
                           A1_21_port);
   U1358 : XOR2X1 port map( A => SUMB_15_9_port, B => CARRYB_15_8_port, Y => 
                           A1_22_port);
   U1359 : XOR2X1 port map( A => SUMB_15_10_port, B => CARRYB_15_9_port, Y => 
                           A1_23_port);
   U1360 : XOR2X1 port map( A => SUMB_15_11_port, B => CARRYB_15_10_port, Y => 
                           A1_24_port);
   U1361 : XOR2X1 port map( A => SUMB_15_12_port, B => CARRYB_15_11_port, Y => 
                           A1_25_port);
   U1362 : XOR2X1 port map( A => SUMB_15_13_port, B => CARRYB_15_12_port, Y => 
                           A1_26_port);
   U1363 : XOR2X1 port map( A => SUMB_15_14_port, B => CARRYB_15_13_port, Y => 
                           A1_27_port);
   U1364 : XOR2X1 port map( A => SUMB_15_15_port, B => CARRYB_15_14_port, Y => 
                           A1_28_port);
   U1365 : XOR2X1 port map( A => ab_1_0_port, B => ab_0_1_port, Y => PRODUCT(1)
                           );
   U1366 : XOR2X1 port map( A => ab_1_1_port, B => ab_0_2_port, Y => 
                           SUMB_1_1_port);
   U1367 : XOR2X1 port map( A => n964, B => ab_0_3_port, Y => SUMB_1_2_port);
   U1368 : XOR2X1 port map( A => ab_1_3_port, B => ab_0_4_port, Y => 
                           SUMB_1_3_port);
   U1369 : XOR2X1 port map( A => ab_0_5_port, B => n525, Y => SUMB_1_4_port);
   U1370 : XOR2X1 port map( A => ab_1_6_port, B => ab_0_7_port, Y => 
                           SUMB_1_6_port);
   U1371 : XOR2X1 port map( A => n439, B => ab_0_8_port, Y => SUMB_1_7_port);
   U1372 : NAND2X1 port map( A => n184, B => ab_0_10_port, Y => n974);
   U1373 : XOR2X1 port map( A => ab_0_11_port, B => ab_1_10_port, Y => 
                           SUMB_1_10_port);
   U1374 : XOR2X1 port map( A => ab_1_12_port, B => ab_0_13_port, Y => 
                           SUMB_1_12_port);
   U1375 : NAND2X1 port map( A => ab_0_13_port, B => ab_1_12_port, Y => n975);
   U1376 : XOR2X1 port map( A => ab_0_14_port, B => ab_1_13_port, Y => 
                           SUMB_1_13_port);
   U1377 : NAND2X1 port map( A => ab_0_14_port, B => ab_1_13_port, Y => n976);
   U1378 : INVX2 port map( A => n976, Y => CARRYB_1_13_port);
   U1379 : XOR2X1 port map( A => ab_1_14_port, B => ab_0_15_port, Y => 
                           SUMB_1_14_port);
   U1380 : INVX2 port map( A => n996, Y => n997);
   U1381 : INVX2 port map( A => n998, Y => n999);
   U1382 : INVX2 port map( A => B(4), Y => n998);
   U1383 : INVX2 port map( A => n1000, Y => n1001);
   U1384 : INVX2 port map( A => B(5), Y => n1000);
   U1385 : INVX1 port map( A => n984, Y => n1044);
   U1386 : INVX1 port map( A => n985, Y => n1043);
   U1387 : INVX4 port map( A => B(2), Y => n994);
   U1388 : INVX8 port map( A => n990, Y => n991);
   U1389 : INVX8 port map( A => n994, Y => n995);
   U1390 : INVX8 port map( A => n1008, Y => n1009);
   U1391 : INVX8 port map( A => n1012, Y => n1013);
   U1392 : INVX8 port map( A => n1014, Y => n1015);
   U1393 : INVX8 port map( A => n1016, Y => n1017);
   U1394 : INVX8 port map( A => n1018, Y => n1019);
   U1395 : INVX8 port map( A => n1024, Y => n1025);
   U1396 : INVX8 port map( A => n1026, Y => n1027);
   U1397 : INVX8 port map( A => n1028, Y => n1029);
   U1398 : INVX8 port map( A => n1030, Y => n1031);
   U1399 : INVX8 port map( A => n1032, Y => n1033);
   U1400 : INVX8 port map( A => n1034, Y => n1035);
   U1401 : INVX8 port map( A => n1036, Y => n1037);
   U1402 : AND2X2 port map( A => n846, B => n1019, Y => ab_1_14_port);
   U1403 : AND2X2 port map( A => n1019, B => n987, Y => ab_0_14_port);
   U1404 : AND2X2 port map( A => n322, B => n1017, Y => ab_1_13_port);
   U1405 : AND2X2 port map( A => n1017, B => n266, Y => ab_0_13_port);
   U1406 : AND2X2 port map( A => n511, B => n1015, Y => ab_1_12_port);
   U1407 : AND2X2 port map( A => n322, B => n1013, Y => ab_1_11_port);
   U1408 : AND2X2 port map( A => n1013, B => n987, Y => ab_0_11_port);
   U1409 : AND2X2 port map( A => n511, B => B(10), Y => ab_1_10_port);
   U1410 : AND2X2 port map( A => n266, B => B(10), Y => ab_0_10_port);
   U1411 : AND2X2 port map( A => n266, B => B(9), Y => ab_0_9_port);
   U1412 : AND2X2 port map( A => n1007, B => n514, Y => ab_1_8_port);
   U1413 : AND2X2 port map( A => n266, B => n239, Y => ab_0_8_port);
   U1414 : AND2X2 port map( A => B(7), B => n987, Y => ab_0_7_port);
   U1415 : AND2X2 port map( A => B(6), B => n514, Y => ab_1_6_port);
   U1416 : AND2X2 port map( A => n1001, B => n514, Y => ab_1_5_port);
   U1417 : AND2X2 port map( A => n1001, B => n266, Y => ab_0_5_port);
   U1418 : AND2X2 port map( A => n999, B => n987, Y => ab_0_4_port);
   U1419 : AND2X2 port map( A => n997, B => n514, Y => ab_1_3_port);
   U1420 : AND2X2 port map( A => n997, B => n987, Y => ab_0_3_port);
   U1421 : AND2X2 port map( A => n995, B => n987, Y => ab_0_2_port);
   U1422 : AND2X2 port map( A => n993, B => n987, Y => ab_0_1_port);
   U1423 : AND2X2 port map( A => n991, B => n846, Y => ab_1_0_port);
   U1424 : AND2X2 port map( A => n235, B => n1019, Y => ab_2_14_port);
   U1425 : NOR2X1 port map( A => n846, B => n1049, Y => ab_1_15_port);
   U1426 : AND2X2 port map( A => n236, B => n1017, Y => ab_2_13_port);
   U1427 : AND2X2 port map( A => n235, B => n1015, Y => ab_2_12_port);
   U1428 : AND2X2 port map( A => n236, B => n1013, Y => ab_2_11_port);
   U1429 : AND2X2 port map( A => n235, B => n51, Y => ab_2_10_port);
   U1430 : AND2X2 port map( A => n206, B => B(9), Y => ab_2_9_port);
   U1431 : AND2X2 port map( A => n1023, B => B(6), Y => ab_2_6_port);
   U1432 : AND2X2 port map( A => n236, B => n983, Y => ab_2_3_port);
   U1433 : AND2X2 port map( A => n1023, B => n995, Y => ab_2_2_port);
   U1434 : AND2X2 port map( A => n235, B => n991, Y => ab_2_0_port);
   U1435 : AND2X2 port map( A => n1025, B => n1019, Y => ab_3_14_port);
   U1436 : NOR2X1 port map( A => n235, B => n1049, Y => ab_2_15_port);
   U1437 : AND2X2 port map( A => n1025, B => n1017, Y => ab_3_13_port);
   U1438 : AND2X2 port map( A => n1025, B => n1015, Y => ab_3_12_port);
   U1439 : AND2X2 port map( A => n1025, B => n1013, Y => ab_3_11_port);
   U1440 : AND2X2 port map( A => n1025, B => n51, Y => ab_3_10_port);
   U1441 : AND2X2 port map( A => n1025, B => B(7), Y => ab_3_7_port);
   U1442 : AND2X2 port map( A => n1025, B => n1003, Y => ab_3_6_port);
   U1443 : AND2X2 port map( A => n1025, B => n985, Y => ab_3_5_port);
   U1444 : AND2X2 port map( A => n1025, B => n984, Y => ab_3_4_port);
   U1445 : AND2X2 port map( A => n1025, B => n983, Y => ab_3_3_port);
   U1446 : AND2X2 port map( A => n1025, B => n995, Y => ab_3_2_port);
   U1447 : AND2X2 port map( A => n1025, B => n993, Y => ab_3_1_port);
   U1448 : AND2X2 port map( A => n396, B => n991, Y => ab_3_0_port);
   U1449 : AND2X2 port map( A => n1027, B => n1019, Y => ab_4_14_port);
   U1450 : NOR2X1 port map( A => n396, B => n1049, Y => ab_3_15_port);
   U1451 : AND2X2 port map( A => n1027, B => n1017, Y => ab_4_13_port);
   U1452 : AND2X2 port map( A => n1027, B => n1015, Y => ab_4_12_port);
   U1453 : AND2X2 port map( A => n1027, B => n1013, Y => ab_4_11_port);
   U1454 : AND2X2 port map( A => n1027, B => n1011, Y => ab_4_10_port);
   U1455 : AND2X2 port map( A => n1027, B => n1009, Y => ab_4_9_port);
   U1456 : AND2X2 port map( A => n1027, B => n1007, Y => ab_4_8_port);
   U1457 : AND2X2 port map( A => n1027, B => n1005, Y => ab_4_7_port);
   U1458 : AND2X2 port map( A => n1027, B => n1003, Y => ab_4_6_port);
   U1459 : AND2X2 port map( A => n1027, B => n985, Y => ab_4_5_port);
   U1460 : AND2X2 port map( A => n1027, B => n984, Y => ab_4_4_port);
   U1461 : AND2X2 port map( A => n1027, B => n983, Y => ab_4_3_port);
   U1462 : AND2X2 port map( A => n1027, B => n995, Y => ab_4_2_port);
   U1463 : AND2X2 port map( A => n1027, B => n993, Y => ab_4_1_port);
   U1464 : AND2X2 port map( A => n1027, B => n991, Y => ab_4_0_port);
   U1465 : AND2X2 port map( A => n1029, B => n1019, Y => ab_5_14_port);
   U1466 : NOR2X1 port map( A => n1027, B => n1049, Y => ab_4_15_port);
   U1467 : AND2X2 port map( A => n1029, B => n1017, Y => ab_5_13_port);
   U1468 : AND2X2 port map( A => n1029, B => n1015, Y => ab_5_12_port);
   U1469 : AND2X2 port map( A => n1029, B => n1013, Y => ab_5_11_port);
   U1470 : AND2X2 port map( A => n1029, B => n1011, Y => ab_5_10_port);
   U1471 : AND2X2 port map( A => n1029, B => n1009, Y => ab_5_9_port);
   U1472 : AND2X2 port map( A => n1029, B => n1007, Y => ab_5_8_port);
   U1473 : AND2X2 port map( A => n1029, B => n1005, Y => ab_5_7_port);
   U1474 : AND2X2 port map( A => n1029, B => n1003, Y => ab_5_6_port);
   U1475 : AND2X2 port map( A => n1029, B => n985, Y => ab_5_5_port);
   U1476 : AND2X2 port map( A => n1029, B => n984, Y => ab_5_4_port);
   U1477 : AND2X2 port map( A => n1029, B => n983, Y => ab_5_3_port);
   U1478 : AND2X2 port map( A => n1029, B => n995, Y => ab_5_2_port);
   U1479 : AND2X2 port map( A => n1029, B => n993, Y => ab_5_1_port);
   U1480 : AND2X2 port map( A => n1029, B => n991, Y => ab_5_0_port);
   U1481 : AND2X2 port map( A => n1031, B => n1019, Y => ab_6_14_port);
   U1482 : NOR2X1 port map( A => n1029, B => n1049, Y => ab_5_15_port);
   U1483 : AND2X2 port map( A => n1031, B => n1017, Y => ab_6_13_port);
   U1484 : AND2X2 port map( A => n1031, B => n1015, Y => ab_6_12_port);
   U1485 : AND2X2 port map( A => n1031, B => n1013, Y => ab_6_11_port);
   U1486 : AND2X2 port map( A => n1031, B => n1011, Y => ab_6_10_port);
   U1487 : AND2X2 port map( A => n1031, B => n1009, Y => ab_6_9_port);
   U1488 : AND2X2 port map( A => n1031, B => n1007, Y => ab_6_8_port);
   U1489 : AND2X2 port map( A => n1031, B => n1005, Y => ab_6_7_port);
   U1490 : AND2X2 port map( A => n1031, B => n1003, Y => ab_6_6_port);
   U1491 : AND2X2 port map( A => n1031, B => n985, Y => ab_6_5_port);
   U1492 : AND2X2 port map( A => n1031, B => n984, Y => ab_6_4_port);
   U1493 : AND2X2 port map( A => n1031, B => n983, Y => ab_6_3_port);
   U1494 : AND2X2 port map( A => n1031, B => n995, Y => ab_6_2_port);
   U1495 : AND2X2 port map( A => n1031, B => n993, Y => ab_6_1_port);
   U1496 : AND2X2 port map( A => n1031, B => n991, Y => ab_6_0_port);
   U1497 : AND2X2 port map( A => n1033, B => n1019, Y => ab_7_14_port);
   U1498 : NOR2X1 port map( A => n1031, B => n1049, Y => ab_6_15_port);
   U1499 : AND2X2 port map( A => n1033, B => n1017, Y => ab_7_13_port);
   U1500 : AND2X2 port map( A => n1033, B => n1015, Y => ab_7_12_port);
   U1501 : AND2X2 port map( A => n1033, B => n1013, Y => ab_7_11_port);
   U1502 : AND2X2 port map( A => n1033, B => n1011, Y => ab_7_10_port);
   U1503 : AND2X2 port map( A => n1033, B => n1009, Y => ab_7_9_port);
   U1504 : AND2X2 port map( A => n1033, B => n132, Y => ab_7_8_port);
   U1505 : AND2X2 port map( A => n1033, B => n1005, Y => ab_7_7_port);
   U1506 : AND2X2 port map( A => n1033, B => n1003, Y => ab_7_6_port);
   U1507 : AND2X2 port map( A => n1033, B => n985, Y => ab_7_5_port);
   U1508 : AND2X2 port map( A => n1033, B => n984, Y => ab_7_4_port);
   U1509 : AND2X2 port map( A => n1033, B => n983, Y => ab_7_3_port);
   U1510 : AND2X2 port map( A => n1033, B => n995, Y => ab_7_2_port);
   U1511 : AND2X2 port map( A => n1033, B => n993, Y => ab_7_1_port);
   U1512 : AND2X2 port map( A => n1033, B => n991, Y => ab_7_0_port);
   U1513 : AND2X2 port map( A => n1035, B => n1019, Y => ab_8_14_port);
   U1514 : NOR2X1 port map( A => n1033, B => n1049, Y => ab_7_15_port);
   U1515 : AND2X2 port map( A => n1035, B => n1017, Y => ab_8_13_port);
   U1516 : AND2X2 port map( A => n1035, B => n1015, Y => ab_8_12_port);
   U1517 : AND2X2 port map( A => n1035, B => n1013, Y => ab_8_11_port);
   U1518 : AND2X2 port map( A => n1035, B => n1011, Y => ab_8_10_port);
   U1519 : AND2X2 port map( A => n1035, B => n1009, Y => ab_8_9_port);
   U1520 : AND2X2 port map( A => n1035, B => n132, Y => ab_8_8_port);
   U1521 : AND2X2 port map( A => n1035, B => n1005, Y => ab_8_7_port);
   U1522 : AND2X2 port map( A => n1035, B => n1003, Y => ab_8_6_port);
   U1523 : AND2X2 port map( A => n1035, B => n985, Y => ab_8_5_port);
   U1524 : AND2X2 port map( A => n1035, B => n984, Y => ab_8_4_port);
   U1525 : AND2X2 port map( A => n1035, B => n983, Y => ab_8_3_port);
   U1526 : AND2X2 port map( A => n1035, B => n995, Y => ab_8_2_port);
   U1527 : AND2X2 port map( A => n1035, B => n993, Y => ab_8_1_port);
   U1528 : AND2X2 port map( A => n1035, B => n991, Y => ab_8_0_port);
   U1529 : AND2X2 port map( A => n1037, B => n1019, Y => ab_9_14_port);
   U1530 : NOR2X1 port map( A => n1035, B => n1049, Y => ab_8_15_port);
   U1531 : AND2X2 port map( A => n1037, B => n1017, Y => ab_9_13_port);
   U1532 : AND2X2 port map( A => n1037, B => n1015, Y => ab_9_12_port);
   U1533 : AND2X2 port map( A => n1037, B => n1013, Y => ab_9_11_port);
   U1534 : AND2X2 port map( A => n1037, B => n1011, Y => ab_9_10_port);
   U1535 : AND2X2 port map( A => n1037, B => n1009, Y => ab_9_9_port);
   U1536 : AND2X2 port map( A => n1037, B => n132, Y => ab_9_8_port);
   U1537 : AND2X2 port map( A => n1037, B => n1005, Y => ab_9_7_port);
   U1538 : AND2X2 port map( A => n1037, B => n1003, Y => ab_9_6_port);
   U1539 : AND2X2 port map( A => n1037, B => n985, Y => ab_9_5_port);
   U1540 : AND2X2 port map( A => n1037, B => n984, Y => ab_9_4_port);
   U1541 : AND2X2 port map( A => n1037, B => n983, Y => ab_9_3_port);
   U1542 : AND2X2 port map( A => n1037, B => n995, Y => ab_9_2_port);
   U1543 : AND2X2 port map( A => n1037, B => n993, Y => ab_9_1_port);
   U1544 : AND2X2 port map( A => n1037, B => n991, Y => ab_9_0_port);
   U1545 : AND2X2 port map( A => A(10), B => n1019, Y => ab_10_14_port);
   U1546 : NOR2X1 port map( A => n1037, B => n1049, Y => ab_9_15_port);
   U1547 : AND2X2 port map( A => A(10), B => n1017, Y => ab_10_13_port);
   U1548 : AND2X2 port map( A => A(10), B => n1015, Y => ab_10_12_port);
   U1549 : AND2X2 port map( A => A(10), B => n1013, Y => ab_10_11_port);
   U1550 : AND2X2 port map( A => A(10), B => n1011, Y => ab_10_10_port);
   U1551 : AND2X2 port map( A => A(10), B => n1009, Y => ab_10_9_port);
   U1552 : AND2X2 port map( A => A(10), B => n132, Y => ab_10_8_port);
   U1553 : AND2X2 port map( A => A(10), B => n1005, Y => ab_10_7_port);
   U1554 : AND2X2 port map( A => A(10), B => n1003, Y => ab_10_6_port);
   U1555 : AND2X2 port map( A => A(10), B => n985, Y => ab_10_5_port);
   U1556 : AND2X2 port map( A => A(10), B => n984, Y => ab_10_4_port);
   U1557 : AND2X2 port map( A => A(10), B => n983, Y => ab_10_3_port);
   U1558 : AND2X2 port map( A => A(10), B => n995, Y => ab_10_2_port);
   U1559 : AND2X2 port map( A => A(10), B => n993, Y => ab_10_1_port);
   U1560 : AND2X2 port map( A => A(10), B => n991, Y => ab_10_0_port);
   U1561 : AND2X2 port map( A => A(11), B => n1019, Y => ab_11_14_port);
   U1562 : NOR2X1 port map( A => A(10), B => n1049, Y => ab_10_15_port);
   U1563 : AND2X2 port map( A => A(11), B => n1017, Y => ab_11_13_port);
   U1564 : AND2X2 port map( A => A(11), B => n1015, Y => ab_11_12_port);
   U1565 : AND2X2 port map( A => A(11), B => n1013, Y => ab_11_11_port);
   U1566 : AND2X2 port map( A => A(11), B => n1011, Y => ab_11_10_port);
   U1567 : AND2X2 port map( A => A(11), B => n1009, Y => ab_11_9_port);
   U1568 : AND2X2 port map( A => A(11), B => n132, Y => ab_11_8_port);
   U1569 : AND2X2 port map( A => A(11), B => n1005, Y => ab_11_7_port);
   U1570 : AND2X2 port map( A => A(11), B => n1003, Y => ab_11_6_port);
   U1571 : AND2X2 port map( A => A(11), B => n985, Y => ab_11_5_port);
   U1572 : AND2X2 port map( A => A(11), B => n984, Y => ab_11_4_port);
   U1573 : AND2X2 port map( A => A(11), B => n983, Y => ab_11_3_port);
   U1574 : AND2X2 port map( A => A(11), B => n995, Y => ab_11_2_port);
   U1575 : AND2X2 port map( A => A(11), B => n993, Y => ab_11_1_port);
   U1576 : AND2X2 port map( A => A(11), B => n991, Y => ab_11_0_port);
   U1577 : AND2X2 port map( A => A(12), B => n1019, Y => ab_12_14_port);
   U1578 : NOR2X1 port map( A => A(11), B => n1049, Y => ab_11_15_port);
   U1579 : AND2X2 port map( A => A(12), B => n1017, Y => ab_12_13_port);
   U1580 : AND2X2 port map( A => A(12), B => n1015, Y => ab_12_12_port);
   U1581 : AND2X2 port map( A => A(12), B => n1013, Y => ab_12_11_port);
   U1582 : AND2X2 port map( A => A(12), B => n1011, Y => ab_12_10_port);
   U1583 : AND2X2 port map( A => A(12), B => n1009, Y => ab_12_9_port);
   U1584 : AND2X2 port map( A => A(12), B => n132, Y => ab_12_8_port);
   U1585 : AND2X2 port map( A => A(12), B => n1005, Y => ab_12_7_port);
   U1586 : AND2X2 port map( A => A(12), B => n1003, Y => ab_12_6_port);
   U1587 : AND2X2 port map( A => A(12), B => n985, Y => ab_12_5_port);
   U1588 : AND2X2 port map( A => A(12), B => n984, Y => ab_12_4_port);
   U1589 : AND2X2 port map( A => A(12), B => n983, Y => ab_12_3_port);
   U1590 : AND2X2 port map( A => A(12), B => n995, Y => ab_12_2_port);
   U1591 : AND2X2 port map( A => A(12), B => n993, Y => ab_12_1_port);
   U1592 : AND2X2 port map( A => A(12), B => n991, Y => ab_12_0_port);
   U1593 : NOR2X1 port map( A => n1052, B => n1018, Y => ab_13_14_port);
   U1594 : NOR2X1 port map( A => A(12), B => n1049, Y => ab_12_15_port);
   U1595 : NOR2X1 port map( A => n1052, B => n1038, Y => ab_13_13_port);
   U1596 : NOR2X1 port map( A => n1052, B => n1039, Y => ab_13_12_port);
   U1597 : NOR2X1 port map( A => n1052, B => n1040, Y => ab_13_11_port);
   U1598 : NOR2X1 port map( A => n1052, B => n1010, Y => ab_13_10_port);
   U1599 : NOR2X1 port map( A => n1052, B => n1041, Y => ab_13_9_port);
   U1600 : NOR2X1 port map( A => n1052, B => n1042, Y => ab_13_8_port);
   U1601 : NOR2X1 port map( A => n1052, B => n1004, Y => ab_13_7_port);
   U1602 : NOR2X1 port map( A => n1052, B => n1002, Y => ab_13_6_port);
   U1603 : NOR2X1 port map( A => n1052, B => n1043, Y => ab_13_5_port);
   U1604 : NOR2X1 port map( A => n1052, B => n1044, Y => ab_13_4_port);
   U1605 : NOR2X1 port map( A => n1052, B => n996, Y => ab_13_3_port);
   U1606 : INVX2 port map( A => n995, Y => n1045);
   U1607 : NOR2X1 port map( A => n1052, B => n1045, Y => ab_13_2_port);
   U1608 : INVX2 port map( A => n993, Y => n1046);
   U1609 : NOR2X1 port map( A => n1052, B => n1046, Y => ab_13_1_port);
   U1610 : INVX2 port map( A => n991, Y => n1047);
   U1611 : NOR2X1 port map( A => n1052, B => n1047, Y => ab_13_0_port);
   U1612 : NOR2X1 port map( A => n1051, B => n1018, Y => ab_14_14_port);
   U1613 : NOR2X1 port map( A => A(13), B => n1049, Y => ab_13_15_port);
   U1614 : NOR2X1 port map( A => n1051, B => n1038, Y => ab_14_13_port);
   U1615 : NOR2X1 port map( A => n1051, B => n1039, Y => ab_14_12_port);
   U1616 : NOR2X1 port map( A => n1051, B => n1040, Y => ab_14_11_port);
   U1617 : NOR2X1 port map( A => n1051, B => n1010, Y => ab_14_10_port);
   U1618 : NOR2X1 port map( A => n1051, B => n1041, Y => ab_14_9_port);
   U1619 : NOR2X1 port map( A => n1051, B => n1042, Y => ab_14_8_port);
   U1620 : NOR2X1 port map( A => n1051, B => n1004, Y => ab_14_7_port);
   U1621 : NOR2X1 port map( A => n1051, B => n1002, Y => ab_14_6_port);
   U1622 : NOR2X1 port map( A => n1051, B => n1043, Y => ab_14_5_port);
   U1623 : NOR2X1 port map( A => n1051, B => n1044, Y => ab_14_4_port);
   U1624 : NOR2X1 port map( A => n1051, B => n996, Y => ab_14_3_port);
   U1625 : NOR2X1 port map( A => n1051, B => n1045, Y => ab_14_2_port);
   U1626 : NOR2X1 port map( A => n1051, B => n1046, Y => ab_14_1_port);
   U1627 : NOR2X1 port map( A => n1051, B => n1047, Y => ab_14_0_port);
   U1628 : NOR2X1 port map( A => n1050, B => n1049, Y => ab_15_15_port);
   U1629 : NOR2X1 port map( A => A(14), B => n1049, Y => ab_14_15_port);
   U1630 : AND2X2 port map( A => n991, B => n987, Y => PRODUCT(0));
   U1631 : INVX2 port map( A => CARRYB_15_15_port, Y => n1048);
   U1632 : NOR2X1 port map( A => n1009, B => n1050, Y => ab_15_9_port);
   U1633 : NOR2X1 port map( A => n132, B => n1050, Y => ab_15_8_port);
   U1634 : NOR2X1 port map( A => n1005, B => n1050, Y => ab_15_7_port);
   U1635 : NOR2X1 port map( A => n1003, B => n1050, Y => ab_15_6_port);
   U1636 : NOR2X1 port map( A => n985, B => n1050, Y => ab_15_5_port);
   U1637 : NOR2X1 port map( A => n984, B => n1050, Y => ab_15_4_port);
   U1638 : NOR2X1 port map( A => n983, B => n1050, Y => ab_15_3_port);
   U1639 : NOR2X1 port map( A => n995, B => n1050, Y => ab_15_2_port);
   U1640 : NOR2X1 port map( A => n993, B => n1050, Y => ab_15_1_port);
   U1641 : NOR2X1 port map( A => n1019, B => n1050, Y => ab_15_14_port);
   U1642 : NOR2X1 port map( A => n1017, B => n1050, Y => ab_15_13_port);
   U1643 : NOR2X1 port map( A => n1015, B => n1050, Y => ab_15_12_port);
   U1644 : NOR2X1 port map( A => n1013, B => n1050, Y => ab_15_11_port);
   U1645 : NOR2X1 port map( A => n1011, B => n1050, Y => ab_15_10_port);
   U1646 : NOR2X1 port map( A => n991, B => n1050, Y => ab_15_0_port);
   n1053 <= '0';

end SYN_csa;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_add_3 is

   port( A, B : in std_logic_vector (8 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (8 downto 0);  CO : out std_logic);

end Rasterizer_DW01_add_3;

architecture SYN_rpl of Rasterizer_DW01_add_3 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port,
      carry_3_port, carry_2_port, n1, n2 : std_logic;

begin
   
   U1_8 : FAX1 port map( A => A(8), B => B(8), C => carry_8_port, YC => n2, YS 
                           => SUM(8));
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => 
                           carry_8_port, YS => SUM(7));
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n1, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_sub_6 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end Rasterizer_DW01_sub_6;

architecture SYN_rpl of Rasterizer_DW01_sub_6 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9 : 
      std_logic;

begin
   
   U2_7 : FAX1 port map( A => A(7), B => n1, C => carry_7_port, YC => n9, YS =>
                           DIFF(7));
   U2_6 : FAX1 port map( A => A(6), B => n2, C => carry_6_port, YC => 
                           carry_7_port, YS => DIFF(6));
   U2_5 : FAX1 port map( A => A(5), B => n3, C => carry_5_port, YC => 
                           carry_6_port, YS => DIFF(5));
   U2_4 : FAX1 port map( A => A(4), B => n4, C => carry_4_port, YC => 
                           carry_5_port, YS => DIFF(4));
   U2_3 : FAX1 port map( A => A(3), B => n5, C => carry_3_port, YC => 
                           carry_4_port, YS => DIFF(3));
   U2_2 : FAX1 port map( A => A(2), B => n6, C => carry_2_port, YC => 
                           carry_3_port, YS => DIFF(2));
   U2_1 : FAX1 port map( A => A(1), B => n7, C => carry_1_port, YC => 
                           carry_2_port, YS => DIFF(1));
   U1 : OR2X2 port map( A => A(0), B => n8, Y => carry_1_port);
   U2 : XNOR2X1 port map( A => n8, B => A(0), Y => DIFF(0));
   U3 : INVX2 port map( A => B(7), Y => n1);
   U4 : INVX2 port map( A => B(6), Y => n2);
   U5 : INVX2 port map( A => B(5), Y => n3);
   U6 : INVX2 port map( A => B(4), Y => n4);
   U7 : INVX2 port map( A => B(3), Y => n5);
   U8 : INVX2 port map( A => B(2), Y => n6);
   U9 : INVX2 port map( A => B(1), Y => n7);
   U10 : INVX2 port map( A => B(0), Y => n8);

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_sub_5 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end Rasterizer_DW01_sub_5;

architecture SYN_rpl of Rasterizer_DW01_sub_5 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9 : 
      std_logic;

begin
   
   U2_7 : FAX1 port map( A => A(7), B => n1, C => carry_7_port, YC => n9, YS =>
                           DIFF(7));
   U2_6 : FAX1 port map( A => A(6), B => n2, C => carry_6_port, YC => 
                           carry_7_port, YS => DIFF(6));
   U2_5 : FAX1 port map( A => A(5), B => n3, C => carry_5_port, YC => 
                           carry_6_port, YS => DIFF(5));
   U2_4 : FAX1 port map( A => A(4), B => n4, C => carry_4_port, YC => 
                           carry_5_port, YS => DIFF(4));
   U2_3 : FAX1 port map( A => A(3), B => n5, C => carry_3_port, YC => 
                           carry_4_port, YS => DIFF(3));
   U2_2 : FAX1 port map( A => A(2), B => n6, C => carry_2_port, YC => 
                           carry_3_port, YS => DIFF(2));
   U2_1 : FAX1 port map( A => A(1), B => n7, C => carry_1_port, YC => 
                           carry_2_port, YS => DIFF(1));
   U1 : OR2X2 port map( A => A(0), B => n8, Y => carry_1_port);
   U2 : XNOR2X1 port map( A => n8, B => A(0), Y => DIFF(0));
   U3 : INVX2 port map( A => B(7), Y => n1);
   U4 : INVX2 port map( A => B(6), Y => n2);
   U5 : INVX2 port map( A => B(5), Y => n3);
   U6 : INVX2 port map( A => B(4), Y => n4);
   U7 : INVX2 port map( A => B(3), Y => n5);
   U8 : INVX2 port map( A => B(2), Y => n6);
   U9 : INVX2 port map( A => B(1), Y => n7);
   U10 : INVX2 port map( A => B(0), Y => n8);

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_sub_4 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end Rasterizer_DW01_sub_4;

architecture SYN_rpl of Rasterizer_DW01_sub_4 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9 : 
      std_logic;

begin
   
   U2_7 : FAX1 port map( A => A(7), B => n1, C => carry_7_port, YC => n9, YS =>
                           DIFF(7));
   U2_6 : FAX1 port map( A => A(6), B => n2, C => carry_6_port, YC => 
                           carry_7_port, YS => DIFF(6));
   U2_5 : FAX1 port map( A => A(5), B => n3, C => carry_5_port, YC => 
                           carry_6_port, YS => DIFF(5));
   U2_4 : FAX1 port map( A => A(4), B => n4, C => carry_4_port, YC => 
                           carry_5_port, YS => DIFF(4));
   U2_3 : FAX1 port map( A => A(3), B => n5, C => carry_3_port, YC => 
                           carry_4_port, YS => DIFF(3));
   U2_2 : FAX1 port map( A => A(2), B => n6, C => carry_2_port, YC => 
                           carry_3_port, YS => DIFF(2));
   U2_1 : FAX1 port map( A => A(1), B => n7, C => carry_1_port, YC => 
                           carry_2_port, YS => DIFF(1));
   U1 : INVX1 port map( A => B(7), Y => n1);
   U2 : OR2X2 port map( A => A(0), B => n8, Y => carry_1_port);
   U3 : XNOR2X1 port map( A => n8, B => A(0), Y => DIFF(0));
   U4 : INVX2 port map( A => B(6), Y => n2);
   U5 : INVX2 port map( A => B(5), Y => n3);
   U6 : INVX2 port map( A => B(4), Y => n4);
   U7 : INVX2 port map( A => B(3), Y => n5);
   U8 : INVX2 port map( A => B(2), Y => n6);
   U9 : INVX2 port map( A => B(1), Y => n7);
   U10 : INVX2 port map( A => B(0), Y => n8);

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_sub_3 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end Rasterizer_DW01_sub_3;

architecture SYN_rpl of Rasterizer_DW01_sub_3 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9 : 
      std_logic;

begin
   
   U2_7 : FAX1 port map( A => A(7), B => n1, C => carry_7_port, YC => n9, YS =>
                           DIFF(7));
   U2_6 : FAX1 port map( A => A(6), B => n2, C => carry_6_port, YC => 
                           carry_7_port, YS => DIFF(6));
   U2_5 : FAX1 port map( A => A(5), B => n3, C => carry_5_port, YC => 
                           carry_6_port, YS => DIFF(5));
   U2_4 : FAX1 port map( A => A(4), B => n4, C => carry_4_port, YC => 
                           carry_5_port, YS => DIFF(4));
   U2_3 : FAX1 port map( A => A(3), B => n5, C => carry_3_port, YC => 
                           carry_4_port, YS => DIFF(3));
   U2_2 : FAX1 port map( A => A(2), B => n6, C => carry_2_port, YC => 
                           carry_3_port, YS => DIFF(2));
   U2_1 : FAX1 port map( A => A(1), B => n7, C => carry_1_port, YC => 
                           carry_2_port, YS => DIFF(1));
   U1 : OR2X2 port map( A => A(0), B => n8, Y => carry_1_port);
   U2 : XNOR2X1 port map( A => n8, B => A(0), Y => DIFF(0));
   U3 : INVX2 port map( A => B(7), Y => n1);
   U4 : INVX2 port map( A => B(6), Y => n2);
   U5 : INVX2 port map( A => B(5), Y => n3);
   U6 : INVX2 port map( A => B(4), Y => n4);
   U7 : INVX2 port map( A => B(3), Y => n5);
   U8 : INVX2 port map( A => B(2), Y => n6);
   U9 : INVX2 port map( A => B(1), Y => n7);
   U10 : INVX2 port map( A => B(0), Y => n8);

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_inc_2 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end Rasterizer_DW01_inc_2;

architecture SYN_rpl of Rasterizer_DW01_inc_2 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_sub_2 is

   port( A, B : in std_logic_vector (11 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (11 downto 0);  CO : out std_logic);

end Rasterizer_DW01_sub_2;

architecture SYN_rpl of Rasterizer_DW01_sub_2 is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, carry_1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9 : 
      std_logic;

begin
   
   U2_8 : FAX1 port map( A => A(8), B => n9, C => carry_8_port, YC => 
                           carry_9_port, YS => DIFF(8));
   U2_7 : FAX1 port map( A => A(7), B => n8, C => carry_7_port, YC => 
                           carry_8_port, YS => DIFF(7));
   U2_6 : FAX1 port map( A => A(6), B => n7, C => carry_6_port, YC => 
                           carry_7_port, YS => DIFF(6));
   U2_5 : FAX1 port map( A => A(5), B => n6, C => carry_5_port, YC => 
                           carry_6_port, YS => DIFF(5));
   U2_4 : FAX1 port map( A => A(4), B => n5, C => carry_4_port, YC => 
                           carry_5_port, YS => DIFF(4));
   U2_3 : FAX1 port map( A => A(3), B => n4, C => carry_3_port, YC => 
                           carry_4_port, YS => DIFF(3));
   U2_2 : FAX1 port map( A => A(2), B => n3, C => carry_2_port, YC => 
                           carry_3_port, YS => DIFF(2));
   U2_1 : FAX1 port map( A => A(1), B => n2, C => carry_1_port, YC => 
                           carry_2_port, YS => DIFF(1));
   U1 : OR2X2 port map( A => A(10), B => carry_10_port, Y => carry_11_port);
   U2 : XNOR2X1 port map( A => carry_10_port, B => A(10), Y => DIFF(10));
   U3 : XNOR2X1 port map( A => A(11), B => carry_11_port, Y => DIFF(11));
   U4 : OR2X2 port map( A => A(9), B => carry_9_port, Y => carry_10_port);
   U5 : XNOR2X1 port map( A => carry_9_port, B => A(9), Y => DIFF(9));
   U6 : OR2X2 port map( A => A(0), B => n1, Y => carry_1_port);
   U7 : XNOR2X1 port map( A => n1, B => A(0), Y => DIFF(0));
   U8 : INVX2 port map( A => B(0), Y => n1);
   U9 : INVX2 port map( A => B(1), Y => n2);
   U10 : INVX2 port map( A => B(2), Y => n3);
   U11 : INVX2 port map( A => B(3), Y => n4);
   U12 : INVX2 port map( A => B(4), Y => n5);
   U13 : INVX2 port map( A => B(5), Y => n6);
   U14 : INVX2 port map( A => B(6), Y => n7);
   U15 : INVX2 port map( A => B(7), Y => n8);
   U16 : INVX2 port map( A => B(8), Y => n9);

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_inc_1 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end Rasterizer_DW01_inc_1;

architecture SYN_rpl of Rasterizer_DW01_inc_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_add_0 is

   port( A, B : in std_logic_vector (11 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (11 downto 0);  CO : out std_logic);

end Rasterizer_DW01_add_0;

architecture SYN_rpl of Rasterizer_DW01_add_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component FAX1
      port( A, B, C : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port,
      carry_4_port, carry_3_port, carry_2_port, n1, n2, n3 : std_logic;

begin
   
   U1_8 : FAX1 port map( A => A(8), B => B(8), C => carry_8_port, YC => 
                           carry_9_port, YS => SUM(8));
   U1_7 : FAX1 port map( A => A(7), B => B(7), C => carry_7_port, YC => 
                           carry_8_port, YS => SUM(7));
   U1_6 : FAX1 port map( A => A(6), B => B(6), C => carry_6_port, YC => 
                           carry_7_port, YS => SUM(6));
   U1_5 : FAX1 port map( A => A(5), B => B(5), C => carry_5_port, YC => 
                           carry_6_port, YS => SUM(5));
   U1_4 : FAX1 port map( A => A(4), B => B(4), C => carry_4_port, YC => 
                           carry_5_port, YS => SUM(4));
   U1_3 : FAX1 port map( A => A(3), B => B(3), C => carry_3_port, YC => 
                           carry_4_port, YS => SUM(3));
   U1_2 : FAX1 port map( A => A(2), B => B(2), C => carry_2_port, YC => 
                           carry_3_port, YS => SUM(2));
   U1_1 : FAX1 port map( A => A(1), B => B(1), C => n1, YC => carry_2_port, YS 
                           => SUM(1));
   U1 : AND2X2 port map( A => B(0), B => A(0), Y => n1);
   U2 : AND2X2 port map( A => carry_9_port, B => A(9), Y => n2);
   U3 : AND2X2 port map( A => n2, B => A(10), Y => n3);
   U4 : XOR2X1 port map( A => A(11), B => n3, Y => SUM(11));
   U5 : XOR2X1 port map( A => n2, B => A(10), Y => SUM(10));
   U6 : XOR2X1 port map( A => carry_9_port, B => A(9), Y => SUM(9));
   U7 : XOR2X1 port map( A => B(0), B => A(0), Y => SUM(0));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer_DW01_inc_0 is

   port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector (7 
         downto 0));

end Rasterizer_DW01_inc_0;

architecture SYN_rpl of Rasterizer_DW01_inc_0 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port : std_logic;

begin
   
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_7_port, B => A(7), Y => SUM(7));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity gpu_controller_DW01_inc_1 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end gpu_controller_DW01_inc_1;

architecture SYN_rpl of gpu_controller_DW01_inc_1 is

   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HAX1 port map( A => A(14), B => carry_14_port, YC => carry_15_port
                           , YS => SUM(14));
   U1_1_13 : HAX1 port map( A => A(13), B => carry_13_port, YC => carry_14_port
                           , YS => SUM(13));
   U1_1_12 : HAX1 port map( A => A(12), B => carry_12_port, YC => carry_13_port
                           , YS => SUM(12));
   U1_1_11 : HAX1 port map( A => A(11), B => carry_11_port, YC => carry_12_port
                           , YS => SUM(11));
   U1_1_10 : HAX1 port map( A => A(10), B => carry_10_port, YC => carry_11_port
                           , YS => SUM(10));
   U1_1_9 : HAX1 port map( A => A(9), B => carry_9_port, YC => carry_10_port, 
                           YS => SUM(9));
   U1_1_8 : HAX1 port map( A => A(8), B => carry_8_port, YC => carry_9_port, YS
                           => SUM(8));
   U1_1_7 : HAX1 port map( A => A(7), B => carry_7_port, YC => carry_8_port, YS
                           => SUM(7));
   U1_1_6 : HAX1 port map( A => A(6), B => carry_6_port, YC => carry_7_port, YS
                           => SUM(6));
   U1_1_5 : HAX1 port map( A => A(5), B => carry_5_port, YC => carry_6_port, YS
                           => SUM(5));
   U1_1_4 : HAX1 port map( A => A(4), B => carry_4_port, YC => carry_5_port, YS
                           => SUM(4));
   U1_1_3 : HAX1 port map( A => A(3), B => carry_3_port, YC => carry_4_port, YS
                           => SUM(3));
   U1_1_2 : HAX1 port map( A => A(2), B => carry_2_port, YC => carry_3_port, YS
                           => SUM(2));
   U1_1_1 : HAX1 port map( A => A(1), B => A(0), YC => carry_2_port, YS => 
                           SUM(1));
   U1 : INVX2 port map( A => A(0), Y => SUM(0));
   U2 : XOR2X1 port map( A => carry_15_port, B => A(15), Y => SUM(15));

end SYN_rpl;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity gpu_controller is

   port( databus : inout std_logic_vector (15 downto 0);  strb_in, clk, rst_n :
         in std_logic;  gpu_done : out std_logic;  ram_in_use, rast_done : in 
         std_logic;  init_rast : out std_logic;  rast_addr : in 
         std_logic_vector (15 downto 0);  rast_strb : in std_logic;  rast_index
         : in std_logic_vector (3 downto 0);  math_done : in std_logic;  
         init_math, strb_matrix, strb_cor : out std_logic;  err : in std_logic;
         addr_out : out std_logic_vector (14 downto 0);  re_out, we_out : out 
         std_logic;  databus_out, opp : out std_logic_vector (15 downto 0));

end gpu_controller;

architecture SYN_struct of gpu_controller is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component TBUFX1
      port( A, EN : in std_logic;  Y : out std_logic);
   end component;
   
   component HAX1
      port( A, B : in std_logic;  YC, YS : out std_logic);
   end component;
   
   component gpu_controller_DW01_inc_1
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal opp_15_port, opp_14_port, opp_13_port, opp_12_port, opp_11_port, 
      opp_10_port, opp_9_port, opp_8_port, opp_7_port, opp_6_port, opp_5_port, 
      opp_4_port, opp_3_port, opp_2_port, opp_1_port, opp_0_port, re, we, 
      state_3_port, state_2_port, state_1_port, state_0_port, addr_15_port, 
      addr_14_port, addr_13_port, addr_12_port, addr_11_port, addr_10_port, 
      addr_9_port, addr_8_port, addr_7_port, addr_6_port, addr_5_port, 
      addr_4_port, addr_3_port, addr_2_port, addr_1_port, addr_0_port, tem, 
      tem2, counter_4_port, counter_3_port, counter_2_port, counter_1_port, 
      counter_0_port, data_reg_15_port, data_reg_14_port, data_reg_13_port, 
      data_reg_12_port, data_reg_11_port, data_reg_10_port, data_reg_9_port, 
      data_reg_8_port, data_reg_7_port, data_reg_6_port, data_reg_5_port, 
      data_reg_4_port, data_reg_3_port, data_reg_2_port, data_reg_1_port, 
      data_reg_0_port, nextre, N297, N298, N299, N300, N301, N302, N303, N304, 
      N305, N306, N307, N308, N309, N310, N311, N312, N314, N315, N316, N317, 
      n1, n2, n3, n7, n8, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
      , n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, 
      n38, n39, n40, n41, n42, n43, n44, n45, n46, n48, n49, n51, n52, n53, n54
      , n59, n61, n63, n65, n67, n68, n69, n73, n74, n75, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86, n87, n88, n90, n91, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n104, n105, n107, n108, n109, n110, n111, 
      n112, n114, n115, n116, n117, n119, n120, n122, n123, n124, n126, n127, 
      n128, n129, n130, n132, n133, n134, n135, n137, n138, n140, n141, n142, 
      n143, n144, n146, n147, n149, n150, n151, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n165, n166, n167, n169, n170, n171, n172, 
      n173, n174, n176, n177, n178, n180, n182, n183, n184, n185, n186, n187, 
      n189, n190, n193, n194, n195, n196, n197, n198, n199, n200, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n293, n294, n295, 
      n296, n297_port, n298_port, n300_port, n312_port, n314_port, n324, n326, 
      n328, n329, n330, n331, add_213_carry_2_port, add_213_carry_3_port, 
      add_213_carry_4_port, n4, n5, n6, n9, n10, n11, n12, n47, n50, n55, n56, 
      n57, n58, n60, n62, n64, n66, n70, n71, n72, n76, n89, n92, n103, n106, 
      n113, n118, n121, n125, n131, n136, n139, n145, n148, n152, n153, n164, 
      n168, n175, n179, n181, n188, n191, n192, n201, n211, n212, n213, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n275, n292, n299_port, n301_port, n302_port, n303_port, n304_port, 
      n305_port, n306_port, n307_port, n308_port, n309_port, n310_port, 
      n311_port, n313, n315_port, n316_port, n317_port, n318, n319, n320, n321,
      n322, n323, n325, n327, n332, n333 : std_logic;

begin
   databus_out <= ( databus(15), databus(14), databus(13), databus(12), 
      databus(11), databus(10), databus(9), databus(8), databus(7), databus(6),
      databus(5), databus(4), databus(3), databus(2), databus(1), databus(0) );
   opp <= ( opp_15_port, opp_14_port, opp_13_port, opp_12_port, opp_11_port, 
      opp_10_port, opp_9_port, opp_8_port, opp_7_port, opp_6_port, opp_5_port, 
      opp_4_port, opp_3_port, opp_2_port, opp_1_port, opp_0_port );
   
   tem_reg : DFFSR port map( D => strb_in, CLK => clk, R => rst_n, S => n273, Q
                           => tem);
   tem2_reg : DFFSR port map( D => tem, CLK => clk, R => rst_n, S => n272, Q =>
                           tem2);
   we_reg : DFFSR port map( D => n274, CLK => clk, R => rst_n, S => n271, Q => 
                           we);
   opcode_reg_15_inst : DFFSR port map( D => n125, CLK => clk, R => rst_n, S =>
                           n270, Q => opp_15_port);
   state_reg_3_inst : DFFSR port map( D => n331, CLK => clk, R => rst_n, S => 
                           n269, Q => state_3_port);
   counter_reg_4_inst : DFFSR port map( D => n293, CLK => clk, R => rst_n, S =>
                           n268, Q => counter_4_port);
   state_reg_2_inst : DFFSR port map( D => n330, CLK => clk, R => rst_n, S => 
                           n267, Q => state_2_port);
   state_reg_0_inst : DFFSR port map( D => n328, CLK => clk, R => rst_n, S => 
                           n266, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => n329, CLK => clk, R => rst_n, S => 
                           n265, Q => state_1_port);
   data_reg_reg_0_inst : DFFPOSX1 port map( D => n103, CLK => clk, Q => 
                           data_reg_0_port);
   data_reg_reg_1_inst : DFFPOSX1 port map( D => n70, CLK => clk, Q => 
                           data_reg_1_port);
   data_reg_reg_2_inst : DFFPOSX1 port map( D => n136, CLK => clk, Q => 
                           data_reg_2_port);
   data_reg_reg_3_inst : DFFPOSX1 port map( D => n66, CLK => clk, Q => 
                           data_reg_3_port);
   data_reg_reg_4_inst : DFFPOSX1 port map( D => n145, CLK => clk, Q => 
                           data_reg_4_port);
   data_reg_reg_5_inst : DFFPOSX1 port map( D => n62, CLK => clk, Q => 
                           data_reg_5_port);
   data_reg_reg_6_inst : DFFPOSX1 port map( D => n148, CLK => clk, Q => 
                           data_reg_6_port);
   data_reg_reg_7_inst : DFFPOSX1 port map( D => n58, CLK => clk, Q => 
                           data_reg_7_port);
   data_reg_reg_8_inst : DFFPOSX1 port map( D => n153, CLK => clk, Q => 
                           data_reg_8_port);
   data_reg_reg_9_inst : DFFPOSX1 port map( D => n57, CLK => clk, Q => 
                           data_reg_9_port);
   data_reg_reg_10_inst : DFFPOSX1 port map( D => n92, CLK => clk, Q => 
                           data_reg_10_port);
   data_reg_reg_11_inst : DFFPOSX1 port map( D => n113, CLK => clk, Q => 
                           data_reg_11_port);
   data_reg_reg_12_inst : DFFPOSX1 port map( D => n76, CLK => clk, Q => 
                           data_reg_12_port);
   data_reg_reg_13_inst : DFFPOSX1 port map( D => n118, CLK => clk, Q => 
                           data_reg_13_port);
   data_reg_reg_14_inst : DFFPOSX1 port map( D => n71, CLK => clk, Q => 
                           data_reg_14_port);
   data_reg_reg_15_inst : DFFPOSX1 port map( D => n121, CLK => clk, Q => 
                           data_reg_15_port);
   opcode_reg_0_inst : DFFSR port map( D => n326, CLK => clk, R => rst_n, S => 
                           n264, Q => opp_0_port);
   opcode_reg_1_inst : DFFSR port map( D => n324, CLK => clk, R => rst_n, S => 
                           n263, Q => opp_1_port);
   opcode_reg_2_inst : DFFSR port map( D => n131, CLK => clk, R => rst_n, S => 
                           n262, Q => opp_2_port);
   opcode_reg_3_inst : DFFSR port map( D => n64, CLK => clk, R => rst_n, S => 
                           n261, Q => opp_3_port);
   opcode_reg_4_inst : DFFSR port map( D => n139, CLK => clk, R => rst_n, S => 
                           n260, Q => opp_4_port);
   opcode_reg_5_inst : DFFSR port map( D => n60, CLK => clk, R => rst_n, S => 
                           n259, Q => opp_5_port);
   opcode_reg_6_inst : DFFSR port map( D => n314_port, CLK => clk, R => rst_n, 
                           S => n258, Q => opp_6_port);
   opcode_reg_7_inst : DFFSR port map( D => n312_port, CLK => clk, R => rst_n, 
                           S => n257, Q => opp_7_port);
   opcode_reg_8_inst : DFFSR port map( D => n152, CLK => clk, R => rst_n, S => 
                           n256, Q => opp_8_port);
   opcode_reg_9_inst : DFFSR port map( D => n56, CLK => clk, R => rst_n, S => 
                           n255, Q => opp_9_port);
   opcode_reg_10_inst : DFFSR port map( D => n89, CLK => clk, R => rst_n, S => 
                           n254, Q => opp_10_port);
   opcode_reg_11_inst : DFFSR port map( D => n106, CLK => clk, R => rst_n, S =>
                           n253, Q => opp_11_port);
   opcode_reg_12_inst : DFFSR port map( D => n72, CLK => clk, R => rst_n, S => 
                           n252, Q => opp_12_port);
   opcode_reg_13_inst : DFFSR port map( D => n300_port, CLK => clk, R => rst_n,
                           S => n251, Q => opp_13_port);
   opcode_reg_14_inst : DFFSR port map( D => n298_port, CLK => clk, R => rst_n,
                           S => n250, Q => opp_14_port);
   counter_reg_3_inst : DFFSR port map( D => n294, CLK => clk, R => rst_n, S =>
                           n249, Q => counter_3_port);
   counter_reg_0_inst : DFFSR port map( D => n297_port, CLK => clk, R => rst_n,
                           S => n248, Q => counter_0_port);
   counter_reg_1_inst : DFFSR port map( D => n296, CLK => clk, R => rst_n, S =>
                           n247, Q => counter_1_port);
   counter_reg_2_inst : DFFSR port map( D => n295, CLK => clk, R => rst_n, S =>
                           n246, Q => counter_2_port);
   addr_reg_15_inst : DFFSR port map( D => n276, CLK => clk, R => rst_n, S => 
                           n245, Q => addr_15_port);
   addr_reg_0_inst : DFFSR port map( D => n291, CLK => clk, R => rst_n, S => 
                           n244, Q => addr_0_port);
   addr_reg_1_inst : DFFSR port map( D => n290, CLK => clk, R => rst_n, S => 
                           n243, Q => addr_1_port);
   addr_reg_2_inst : DFFSR port map( D => n289, CLK => clk, R => rst_n, S => 
                           n242, Q => addr_2_port);
   addr_reg_3_inst : DFFSR port map( D => n288, CLK => clk, R => rst_n, S => 
                           n241, Q => addr_3_port);
   addr_reg_4_inst : DFFSR port map( D => n287, CLK => clk, R => rst_n, S => 
                           n240, Q => addr_4_port);
   addr_reg_5_inst : DFFSR port map( D => n286, CLK => clk, R => rst_n, S => 
                           n239, Q => addr_5_port);
   addr_reg_6_inst : DFFSR port map( D => n285, CLK => clk, R => rst_n, S => 
                           n238, Q => addr_6_port);
   addr_reg_7_inst : DFFSR port map( D => n284, CLK => clk, R => rst_n, S => 
                           n237, Q => addr_7_port);
   addr_reg_8_inst : DFFSR port map( D => n283, CLK => clk, R => rst_n, S => 
                           n236, Q => addr_8_port);
   addr_reg_9_inst : DFFSR port map( D => n282, CLK => clk, R => rst_n, S => 
                           n235, Q => addr_9_port);
   addr_reg_10_inst : DFFSR port map( D => n281, CLK => clk, R => rst_n, S => 
                           n234, Q => addr_10_port);
   addr_reg_11_inst : DFFSR port map( D => n280, CLK => clk, R => rst_n, S => 
                           n233, Q => addr_11_port);
   addr_reg_12_inst : DFFSR port map( D => n279, CLK => clk, R => rst_n, S => 
                           n232, Q => addr_12_port);
   addr_reg_13_inst : DFFSR port map( D => n278, CLK => clk, R => rst_n, S => 
                           n231, Q => addr_13_port);
   addr_reg_14_inst : DFFSR port map( D => n277, CLK => clk, R => rst_n, S => 
                           n230, Q => addr_14_port);
   re_reg : DFFSR port map( D => nextre, CLK => clk, R => rst_n, S => n229, Q 
                           => re);
   U4 : NOR2X1 port map( A => n1, B => n2, Y => strb_matrix);
   U5 : NOR2X1 port map( A => n2, B => n3, Y => strb_cor);
   U6 : OAI21X1 port map( A => n211, B => n322, C => n164, Y => nextre);
   U8 : NAND2X1 port map( A => n7, B => n8, Y => n276);
   U9 : AOI22X1 port map( A => addr_15_port, B => n4, C => N312, D => n179, Y 
                           => n8);
   U10 : AOI22X1 port map( A => rast_addr(15), B => n201, C => databus(15), D 
                           => n212, Y => n7);
   U11 : NAND2X1 port map( A => n13, B => n14, Y => n277);
   U12 : AOI22X1 port map( A => n4, B => addr_14_port, C => N311, D => n179, Y 
                           => n14);
   U13 : AOI22X1 port map( A => rast_addr(14), B => n201, C => databus(14), D 
                           => n212, Y => n13);
   U14 : NAND2X1 port map( A => n15, B => n16, Y => n278);
   U15 : AOI22X1 port map( A => n4, B => addr_13_port, C => N310, D => n179, Y 
                           => n16);
   U16 : AOI22X1 port map( A => rast_addr(13), B => n201, C => databus(13), D 
                           => n212, Y => n15);
   U17 : NAND2X1 port map( A => n17, B => n18, Y => n279);
   U18 : AOI22X1 port map( A => n4, B => addr_12_port, C => N309, D => n179, Y 
                           => n18);
   U19 : AOI22X1 port map( A => rast_addr(12), B => n201, C => databus(12), D 
                           => n212, Y => n17);
   U20 : NAND2X1 port map( A => n19, B => n20, Y => n280);
   U21 : AOI22X1 port map( A => n4, B => addr_11_port, C => N308, D => n179, Y 
                           => n20);
   U22 : AOI22X1 port map( A => rast_addr(11), B => n201, C => databus(11), D 
                           => n212, Y => n19);
   U23 : NAND2X1 port map( A => n21, B => n22, Y => n281);
   U24 : AOI22X1 port map( A => n4, B => addr_10_port, C => N307, D => n179, Y 
                           => n22);
   U25 : AOI22X1 port map( A => rast_addr(10), B => n201, C => databus(10), D 
                           => n212, Y => n21);
   U26 : NAND2X1 port map( A => n23, B => n24, Y => n282);
   U27 : AOI22X1 port map( A => n4, B => addr_9_port, C => N306, D => n179, Y 
                           => n24);
   U28 : AOI22X1 port map( A => rast_addr(9), B => n201, C => databus(9), D => 
                           n212, Y => n23);
   U29 : NAND2X1 port map( A => n25, B => n26, Y => n283);
   U30 : AOI22X1 port map( A => n4, B => addr_8_port, C => N305, D => n179, Y 
                           => n26);
   U31 : AOI22X1 port map( A => rast_addr(8), B => n201, C => databus(8), D => 
                           n212, Y => n25);
   U32 : NAND2X1 port map( A => n27, B => n28, Y => n284);
   U33 : AOI22X1 port map( A => n4, B => addr_7_port, C => N304, D => n179, Y 
                           => n28);
   U34 : AOI22X1 port map( A => rast_addr(7), B => n201, C => databus(7), D => 
                           n212, Y => n27);
   U35 : NAND2X1 port map( A => n29, B => n30, Y => n285);
   U36 : AOI22X1 port map( A => n4, B => addr_6_port, C => N303, D => n179, Y 
                           => n30);
   U37 : AOI22X1 port map( A => rast_addr(6), B => n201, C => databus(6), D => 
                           n212, Y => n29);
   U38 : NAND2X1 port map( A => n31, B => n32, Y => n286);
   U39 : AOI22X1 port map( A => n4, B => addr_5_port, C => N302, D => n179, Y 
                           => n32);
   U40 : AOI22X1 port map( A => rast_addr(5), B => n201, C => databus(5), D => 
                           n212, Y => n31);
   U41 : NAND2X1 port map( A => n33, B => n34, Y => n287);
   U42 : AOI22X1 port map( A => n4, B => addr_4_port, C => N301, D => n179, Y 
                           => n34);
   U43 : AOI22X1 port map( A => rast_addr(4), B => n201, C => databus(4), D => 
                           n212, Y => n33);
   U44 : NAND2X1 port map( A => n35, B => n36, Y => n288);
   U45 : AOI22X1 port map( A => n4, B => addr_3_port, C => N300, D => n179, Y 
                           => n36);
   U46 : AOI22X1 port map( A => rast_addr(3), B => n201, C => databus(3), D => 
                           n212, Y => n35);
   U47 : NAND2X1 port map( A => n37, B => n38, Y => n289);
   U48 : AOI22X1 port map( A => n4, B => addr_2_port, C => N299, D => n179, Y 
                           => n38);
   U49 : AOI22X1 port map( A => rast_addr(2), B => n201, C => databus(2), D => 
                           n212, Y => n37);
   U50 : NAND2X1 port map( A => n39, B => n40, Y => n290);
   U51 : AOI22X1 port map( A => n4, B => addr_1_port, C => N298, D => n179, Y 
                           => n40);
   U52 : AOI22X1 port map( A => rast_addr(1), B => n201, C => databus(1), D => 
                           n212, Y => n39);
   U53 : NAND2X1 port map( A => n41, B => n42, Y => n291);
   U54 : AOI22X1 port map( A => n4, B => addr_0_port, C => N297, D => n179, Y 
                           => n42);
   U56 : NAND3X1 port map( A => n45, B => n46, C => n192, Y => n44);
   U58 : NAND3X1 port map( A => n49, B => n213, C => n51, Y => n43);
   U59 : AOI22X1 port map( A => rast_addr(0), B => n201, C => databus(0), D => 
                           n212, Y => n41);
   U63 : AOI22X1 port map( A => databus(15), B => n11, C => n5, D => 
                           data_reg_15_port, Y => n54);
   U64 : OAI21X1 port map( A => n188, B => n217, C => n59, Y => n293);
   U65 : NAND2X1 port map( A => N317, B => n179, Y => n59);
   U66 : OAI21X1 port map( A => n188, B => n299_port, C => n61, Y => n294);
   U67 : NAND2X1 port map( A => N316, B => n179, Y => n61);
   U68 : OAI21X1 port map( A => n188, B => n303_port, C => n63, Y => n295);
   U69 : NAND2X1 port map( A => N315, B => n179, Y => n63);
   U70 : OAI21X1 port map( A => n188, B => n302_port, C => n65, Y => n296);
   U71 : NAND2X1 port map( A => N314, B => n179, Y => n65);
   U72 : OAI21X1 port map( A => n188, B => n301_port, C => n67, Y => n297_port)
                           ;
   U73 : NAND2X1 port map( A => n301_port, B => n179, Y => n67);
   U75 : NAND3X1 port map( A => n69, B => n213, C => n191, Y => n68);
   U77 : OAI22X1 port map( A => n9, B => n292, C => n73, D => n10, Y => 
                           n298_port);
   U80 : AOI22X1 port map( A => databus(14), B => n11, C => n5, D => 
                           data_reg_14_port, Y => n75);
   U81 : OAI22X1 port map( A => n9, B => n275, C => n77, D => n10, Y => 
                           n300_port);
   U84 : AOI22X1 port map( A => databus(13), B => n11, C => n5, D => 
                           data_reg_13_port, Y => n78);
   U86 : AOI22X1 port map( A => n10, B => opp_12_port, C => databus(12), D => 
                           n9, Y => n79);
   U88 : AOI22X1 port map( A => databus(12), B => n11, C => n5, D => 
                           data_reg_12_port, Y => n80);
   U90 : AOI22X1 port map( A => n74, B => opp_11_port, C => databus(11), D => 
                           n9, Y => n81);
   U92 : AOI22X1 port map( A => databus(11), B => n11, C => n5, D => 
                           data_reg_11_port, Y => n82);
   U94 : AOI22X1 port map( A => n74, B => opp_10_port, C => databus(10), D => 
                           n9, Y => n83);
   U96 : AOI22X1 port map( A => databus(10), B => n11, C => n5, D => 
                           data_reg_10_port, Y => n84);
   U98 : AOI22X1 port map( A => n74, B => opp_9_port, C => databus(9), D => n9,
                           Y => n85);
   U100 : AOI22X1 port map( A => databus(9), B => n11, C => n5, D => 
                           data_reg_9_port, Y => n86);
   U102 : AOI22X1 port map( A => n74, B => opp_8_port, C => databus(8), D => n9
                           , Y => n87);
   U104 : AOI22X1 port map( A => databus(8), B => n11, C => n5, D => 
                           data_reg_8_port, Y => n88);
   U105 : OAI22X1 port map( A => n9, B => n227, C => n90, D => n10, Y => 
                           n312_port);
   U108 : AOI22X1 port map( A => databus(7), B => n11, C => n5, D => 
                           data_reg_7_port, Y => n91);
   U109 : OAI22X1 port map( A => n9, B => n226, C => n93, D => n10, Y => 
                           n314_port);
   U112 : AOI22X1 port map( A => databus(6), B => n11, C => n5, D => 
                           data_reg_6_port, Y => n94);
   U114 : AOI22X1 port map( A => n74, B => opp_5_port, C => databus(5), D => n9
                           , Y => n95);
   U116 : AOI22X1 port map( A => databus(5), B => n11, C => n5, D => 
                           data_reg_5_port, Y => n96);
   U118 : AOI22X1 port map( A => n74, B => opp_4_port, C => databus(4), D => n9
                           , Y => n97);
   U120 : AOI22X1 port map( A => databus(4), B => n11, C => n5, D => 
                           data_reg_4_port, Y => n98);
   U122 : AOI22X1 port map( A => n74, B => opp_3_port, C => databus(3), D => n9
                           , Y => n99);
   U124 : AOI22X1 port map( A => databus(3), B => n11, C => n5, D => 
                           data_reg_3_port, Y => n100);
   U126 : AOI22X1 port map( A => n74, B => opp_2_port, C => databus(2), D => n9
                           , Y => n101);
   U128 : AOI22X1 port map( A => databus(2), B => n11, C => n5, D => 
                           data_reg_2_port, Y => n102);
   U129 : OAI22X1 port map( A => n9, B => n224, C => n104, D => n10, Y => n324)
                           ;
   U132 : AOI22X1 port map( A => databus(1), B => n11, C => n5, D => 
                           data_reg_1_port, Y => n105);
   U133 : OAI22X1 port map( A => n9, B => n223, C => n107, D => n10, Y => n326)
                           ;
   U136 : AOI22X1 port map( A => databus(0), B => n11, C => n5, D => 
                           data_reg_0_port, Y => n108);
   U139 : NAND3X1 port map( A => n191, B => n69, C => rst_n, Y => n110);
   U140 : NAND3X1 port map( A => n46, B => n2, C => n111, Y => n109);
   U141 : OAI21X1 port map( A => n112, B => n221, C => n114, Y => n328);
   U142 : OAI21X1 port map( A => n115, B => n116, C => n112, Y => n114);
   U143 : OAI21X1 port map( A => n117, B => n46, C => n181, Y => n116);
   U145 : NAND2X1 port map( A => n120, B => n111, Y => n115);
   U146 : OAI21X1 port map( A => n112, B => n222, C => n122, Y => n329);
   U147 : OAI21X1 port map( A => n123, B => n124, C => n112, Y => n122);
   U148 : NAND2X1 port map( A => n45, B => n211, Y => n124);
   U149 : NOR2X1 port map( A => n216, B => n126, Y => n45);
   U150 : OAI21X1 port map( A => n127, B => n128, C => n129, Y => n126);
   U152 : NAND2X1 port map( A => n130, B => n218, Y => n69);
   U153 : NAND3X1 port map( A => n132, B => n133, C => n134, Y => n330);
   U154 : NOR2X1 port map( A => n123, B => n135, Y => n134);
   U155 : OAI21X1 port map( A => n112, B => n220, C => n120, Y => n135);
   U157 : NAND3X1 port map( A => counter_2_port, B => counter_1_port, C => n215
                           , Y => n138);
   U159 : NAND3X1 port map( A => n299_port, B => n217, C => n140, Y => n137);
   U160 : NOR2X1 port map( A => counter_0_port, B => n3, Y => n140);
   U162 : OAI21X1 port map( A => err, B => n141, C => n142, Y => n123);
   U164 : AOI21X1 port map( A => n144, B => n164, C => n12, Y => n331);
   U166 : NOR2X1 port map( A => n146, B => n147, Y => n112);
   U167 : OAI22X1 port map( A => n211, B => rast_strb, C => n129, D => n47, Y 
                           => n147);
   U169 : OAI22X1 port map( A => n133, B => n333, C => n141, D => math_done, Y 
                           => n146);
   U171 : OAI21X1 port map( A => n49, B => n151, C => n51, Y => n150);
   U172 : OAI21X1 port map( A => n168, B => n175, C => n154, Y => n151);
   U173 : NAND3X1 port map( A => n301_port, B => n299_port, C => n155, Y => 
                           n154);
   U174 : OAI21X1 port map( A => n156, B => n157, C => n158, Y => n155);
   U175 : NAND3X1 port map( A => counter_2_port, B => counter_1_port, C => n159
                           , Y => n158);
   U176 : NOR2X1 port map( A => counter_4_port, B => n3, Y => n159);
   U177 : NAND2X1 port map( A => counter_4_port, B => n175, Y => n157);
   U178 : NAND2X1 port map( A => n302_port, B => n303_port, Y => n156);
   U184 : NAND3X1 port map( A => n160, B => n224, C => opp_0_port, Y => n1);
   U187 : NAND3X1 port map( A => n160, B => n223, C => opp_1_port, Y => n3);
   U190 : NOR2X1 port map( A => n163, B => n225, Y => n162);
   U192 : NOR3X1 port map( A => opp_4_port, B => opp_5_port, C => opp_3_port, Y
                           => n165);
   U193 : NAND3X1 port map( A => n226, B => n227, C => n166, Y => n163);
   U194 : NOR2X1 port map( A => opp_9_port, B => opp_8_port, Y => n166);
   U197 : NOR2X1 port map( A => n167, B => n228, Y => n161);
   U199 : NOR3X1 port map( A => opp_11_port, B => opp_12_port, C => opp_10_port
                           , Y => n169);
   U200 : NAND3X1 port map( A => n275, B => n292, C => n170, Y => n167);
   U201 : NOR2X1 port map( A => opp_2_port, B => opp_15_port, Y => n170);
   U204 : NOR2X1 port map( A => n274, B => n149, Y => n144);
   U205 : NOR2X1 port map( A => rast_done, B => n53, Y => n149);
   U207 : AOI22X1 port map( A => n10, B => opp_15_port, C => databus(15), D => 
                           n9, Y => n171);
   U209 : NAND3X1 port map( A => n191, B => n46, C => n132, Y => n74);
   U210 : NOR2X1 port map( A => n274, B => n179, Y => n132);
   U212 : NAND3X1 port map( A => n218, B => n222, C => state_3_port, Y => n2);
   U214 : NAND3X1 port map( A => n53, B => n49, C => n173, Y => n172);
   U215 : NOR2X1 port map( A => n48, B => n119, Y => n173);
   U216 : NAND3X1 port map( A => n52, B => n51, C => n129, Y => n119);
   U217 : NAND2X1 port map( A => n174, B => n219, Y => n129);
   U218 : NAND2X1 port map( A => n219, B => state_3_port, Y => n51);
   U219 : NAND2X1 port map( A => n174, B => n218, Y => n52);
   U221 : NAND3X1 port map( A => n141, B => n143, C => n133, Y => n48);
   U222 : NAND3X1 port map( A => state_2_port, B => state_0_port, C => n174, Y 
                           => n133);
   U223 : NAND3X1 port map( A => state_3_port, B => n177, C => state_2_port, Y 
                           => n143);
   U224 : XOR2X1 port map( A => state_1_port, B => state_0_port, Y => n177);
   U225 : NAND3X1 port map( A => n130, B => n221, C => state_2_port, Y => n49);
   U226 : NAND3X1 port map( A => state_2_port, B => n221, C => n174, Y => n53);
   U227 : NOR2X1 port map( A => n222, B => state_3_port, Y => n174);
   U229 : OAI21X1 port map( A => n176, B => n128, C => n111, Y => n274);
   U230 : NAND3X1 port map( A => state_2_port, B => state_3_port, C => n178, Y 
                           => n111);
   U231 : NOR2X1 port map( A => state_1_port, B => state_0_port, Y => n178);
   U232 : NAND2X1 port map( A => state_1_port, B => state_3_port, Y => n128);
   U233 : NAND2X1 port map( A => state_0_port, B => n220, Y => n176);
   U235 : NOR2X1 port map( A => n332, B => n180, Y => init_rast);
   U237 : NAND3X1 port map( A => n130, B => state_0_port, C => state_2_port, Y 
                           => n141);
   U239 : NOR2X1 port map( A => n47, B => n46, Y => gpu_done);
   U240 : NAND2X1 port map( A => n130, B => n219, Y => n46);
   U242 : NAND2X1 port map( A => n220, B => n221, Y => n127);
   U245 : NOR2X1 port map( A => state_3_port, B => state_1_port, Y => n130);
   U247 : NAND2X1 port map( A => tem, B => n50, Y => n117);
   U249 : AOI21X1 port map( A => n182, B => n183, C => data_reg_9_port, Y => 
                           n200);
   U250 : AOI21X1 port map( A => n184, B => n182, C => data_reg_8_port, Y => 
                           n202);
   U251 : AOI21X1 port map( A => n185, B => n186, C => data_reg_7_port, Y => 
                           n203);
   U252 : AOI21X1 port map( A => n187, B => n186, C => data_reg_6_port, Y => 
                           n204);
   U253 : AOI21X1 port map( A => n186, B => n183, C => data_reg_5_port, Y => 
                           n205);
   U254 : AOI21X1 port map( A => n186, B => n184, C => data_reg_4_port, Y => 
                           n206);
   U255 : NOR2X1 port map( A => n323, B => rast_index(3), Y => n186);
   U256 : AOI21X1 port map( A => n189, B => n185, C => data_reg_3_port, Y => 
                           n207);
   U257 : AOI21X1 port map( A => n189, B => n187, C => data_reg_2_port, Y => 
                           n208);
   U258 : AOI21X1 port map( A => n189, B => n183, C => data_reg_1_port, Y => 
                           n209);
   U259 : AOI21X1 port map( A => n190, B => n185, C => data_reg_15_port, Y => 
                           n194);
   U260 : AOI21X1 port map( A => n190, B => n187, C => data_reg_14_port, Y => 
                           n195);
   U261 : AOI21X1 port map( A => n190, B => n183, C => data_reg_13_port, Y => 
                           n196);
   U262 : NOR2X1 port map( A => n327, B => rast_index(1), Y => n183);
   U263 : AOI21X1 port map( A => n190, B => n184, C => data_reg_12_port, Y => 
                           n197);
   U264 : NOR2X1 port map( A => n323, B => n325, Y => n190);
   U266 : AOI21X1 port map( A => n185, B => n182, C => data_reg_11_port, Y => 
                           n198);
   U268 : AOI21X1 port map( A => n187, B => n182, C => data_reg_10_port, Y => 
                           n199);
   U269 : NOR2X1 port map( A => n325, B => rast_index(2), Y => n182);
   U274 : NAND3X1 port map( A => n333, B => n321, C => we, Y => n193);
   U276 : AOI21X1 port map( A => n189, B => n184, C => data_reg_0_port, Y => 
                           n210);
   U277 : NOR2X1 port map( A => rast_index(1), B => rast_index(0), Y => n184);
   U278 : NOR2X1 port map( A => rast_index(3), B => rast_index(2), Y => n189);
   n229 <= '1';
   n230 <= '1';
   n231 <= '1';
   n232 <= '1';
   n233 <= '1';
   n234 <= '1';
   n235 <= '1';
   n236 <= '1';
   n237 <= '1';
   n238 <= '1';
   n239 <= '1';
   n240 <= '1';
   n241 <= '1';
   n242 <= '1';
   n243 <= '1';
   n244 <= '1';
   n245 <= '1';
   n246 <= '1';
   n247 <= '1';
   n248 <= '1';
   n249 <= '1';
   n250 <= '1';
   n251 <= '1';
   n252 <= '1';
   n253 <= '1';
   n254 <= '1';
   n255 <= '1';
   n256 <= '1';
   n257 <= '1';
   n258 <= '1';
   n259 <= '1';
   n260 <= '1';
   n261 <= '1';
   n262 <= '1';
   n263 <= '1';
   n264 <= '1';
   n265 <= '1';
   n266 <= '1';
   n267 <= '1';
   n268 <= '1';
   n269 <= '1';
   n270 <= '1';
   n271 <= '1';
   n272 <= '1';
   n273 <= '1';
   U78 : INVX2 port map( A => databus(14), Y => n73);
   U82 : INVX2 port map( A => databus(13), Y => n77);
   U106 : INVX2 port map( A => databus(7), Y => n90);
   U110 : INVX2 port map( A => databus(6), Y => n93);
   U130 : INVX2 port map( A => databus(1), Y => n104);
   U134 : INVX2 port map( A => databus(0), Y => n107);
   U156 : OR2X2 port map( A => n137, B => n138, Y => n120);
   U163 : AND2X2 port map( A => n143, B => n52, Y => n142);
   U189 : AND2X2 port map( A => n161, B => n162, Y => n160);
   U236 : OR2X2 port map( A => n141, B => err, Y => n180);
   U267 : AND2X2 port map( A => rast_index(1), B => rast_index(0), Y => n185);
   U271 : AND2X2 port map( A => rast_index(1), B => n327, Y => n187);
   add_212 : gpu_controller_DW01_inc_1 port map( A(15) => addr_15_port, A(14) 
                           => addr_14_port, A(13) => addr_13_port, A(12) => 
                           addr_12_port, A(11) => addr_11_port, A(10) => 
                           addr_10_port, A(9) => addr_9_port, A(8) => 
                           addr_8_port, A(7) => addr_7_port, A(6) => 
                           addr_6_port, A(5) => addr_5_port, A(4) => 
                           addr_4_port, A(3) => addr_3_port, A(2) => 
                           addr_2_port, A(1) => addr_1_port, A(0) => 
                           addr_0_port, SUM(15) => N312, SUM(14) => N311, 
                           SUM(13) => N310, SUM(12) => N309, SUM(11) => N308, 
                           SUM(10) => N307, SUM(9) => N306, SUM(8) => N305, 
                           SUM(7) => N304, SUM(6) => N303, SUM(5) => N302, 
                           SUM(4) => N301, SUM(3) => N300, SUM(2) => N299, 
                           SUM(1) => N298, SUM(0) => N297);
   add_213_U1_1_1 : HAX1 port map( A => counter_1_port, B => counter_0_port, YC
                           => add_213_carry_2_port, YS => N314);
   add_213_U1_1_2 : HAX1 port map( A => counter_2_port, B => 
                           add_213_carry_2_port, YC => add_213_carry_3_port, YS
                           => N315);
   add_213_U1_1_3 : HAX1 port map( A => counter_3_port, B => 
                           add_213_carry_3_port, YC => add_213_carry_4_port, YS
                           => N316);
   databus_tri_15_inst : TBUFX1 port map( A => n194, EN => n6, Y => databus(15)
                           );
   databus_tri_14_inst : TBUFX1 port map( A => n195, EN => n6, Y => databus(14)
                           );
   databus_tri_2_inst : TBUFX1 port map( A => n208, EN => n6, Y => databus(2));
   databus_tri_3_inst : TBUFX1 port map( A => n207, EN => n6, Y => databus(3));
   databus_tri_4_inst : TBUFX1 port map( A => n206, EN => n6, Y => databus(4));
   databus_tri_12_inst : TBUFX1 port map( A => n197, EN => n6, Y => databus(12)
                           );
   databus_tri_8_inst : TBUFX1 port map( A => n202, EN => n6, Y => databus(8));
   databus_tri_10_inst : TBUFX1 port map( A => n199, EN => n6, Y => databus(10)
                           );
   databus_tri_11_inst : TBUFX1 port map( A => n198, EN => n6, Y => databus(11)
                           );
   databus_tri_0_inst : TBUFX1 port map( A => n210, EN => n6, Y => databus(0));
   databus_tri_5_inst : TBUFX1 port map( A => n205, EN => n6, Y => databus(5));
   databus_tri_9_inst : TBUFX1 port map( A => n200, EN => n6, Y => databus(9));
   databus_tri_6_inst : TBUFX1 port map( A => n204, EN => n6, Y => databus(6));
   databus_tri_7_inst : TBUFX1 port map( A => n203, EN => n6, Y => databus(7));
   databus_tri_1_inst : TBUFX1 port map( A => n209, EN => n6, Y => databus(1));
   databus_tri_13_inst : TBUFX1 port map( A => n196, EN => n6, Y => databus(13)
                           );
   re_out_tri : TBUFX1 port map( A => n321, EN => n333, Y => re_out);
   we_out_tri : TBUFX1 port map( A => n55, EN => n333, Y => we_out);
   addr_out_tri_1_inst : TBUFX1 port map( A => n305_port, EN => n333, Y => 
                           addr_out(1));
   addr_out_tri_2_inst : TBUFX1 port map( A => n306_port, EN => n333, Y => 
                           addr_out(2));
   addr_out_tri_3_inst : TBUFX1 port map( A => n307_port, EN => n333, Y => 
                           addr_out(3));
   addr_out_tri_4_inst : TBUFX1 port map( A => n308_port, EN => n333, Y => 
                           addr_out(4));
   addr_out_tri_5_inst : TBUFX1 port map( A => n309_port, EN => n333, Y => 
                           addr_out(5));
   addr_out_tri_6_inst : TBUFX1 port map( A => n310_port, EN => n333, Y => 
                           addr_out(6));
   addr_out_tri_7_inst : TBUFX1 port map( A => n311_port, EN => n333, Y => 
                           addr_out(7));
   addr_out_tri_8_inst : TBUFX1 port map( A => n313, EN => n333, Y => 
                           addr_out(8));
   addr_out_tri_9_inst : TBUFX1 port map( A => n315_port, EN => n333, Y => 
                           addr_out(9));
   addr_out_tri_10_inst : TBUFX1 port map( A => n316_port, EN => n333, Y => 
                           addr_out(10));
   addr_out_tri_11_inst : TBUFX1 port map( A => n317_port, EN => n333, Y => 
                           addr_out(11));
   addr_out_tri_12_inst : TBUFX1 port map( A => n318, EN => n333, Y => 
                           addr_out(12));
   addr_out_tri_13_inst : TBUFX1 port map( A => n319, EN => n333, Y => 
                           addr_out(13));
   addr_out_tri_14_inst : TBUFX1 port map( A => n320, EN => n333, Y => 
                           addr_out(14));
   addr_out_tri_0_inst : TBUFX1 port map( A => n304_port, EN => n333, Y => 
                           addr_out(0));
   U3 : OR2X2 port map( A => n43, B => n44, Y => n4);
   U7 : INVX2 port map( A => n9, Y => n10);
   U55 : INVX2 port map( A => n74, Y => n9);
   U57 : INVX2 port map( A => n5, Y => n11);
   U60 : INVX2 port map( A => n52, Y => n212);
   U61 : INVX2 port map( A => n2, Y => n179);
   U62 : OR2X2 port map( A => n109, B => n110, Y => n5);
   U74 : INVX2 port map( A => n53, Y => n201);
   U76 : INVX2 port map( A => n193, Y => n6);
   U79 : INVX2 port map( A => ram_in_use, Y => n333);
   U83 : XOR2X1 port map( A => add_213_carry_4_port, B => counter_4_port, Y => 
                           N317);
   U85 : INVX2 port map( A => n112, Y => n12);
   U87 : INVX2 port map( A => n117, Y => n47);
   U89 : INVX2 port map( A => tem2, Y => n50);
   U91 : INVX2 port map( A => we, Y => n55);
   U93 : INVX2 port map( A => n85, Y => n56);
   U95 : INVX2 port map( A => n86, Y => n57);
   U97 : INVX2 port map( A => n91, Y => n58);
   U99 : INVX2 port map( A => n95, Y => n60);
   U101 : INVX2 port map( A => n96, Y => n62);
   U103 : INVX2 port map( A => n99, Y => n64);
   U107 : INVX2 port map( A => n100, Y => n66);
   U111 : INVX2 port map( A => n105, Y => n70);
   U113 : INVX2 port map( A => n75, Y => n71);
   U115 : INVX2 port map( A => n79, Y => n72);
   U117 : INVX2 port map( A => n80, Y => n76);
   U119 : INVX2 port map( A => n83, Y => n89);
   U121 : INVX2 port map( A => n84, Y => n92);
   U123 : INVX2 port map( A => n108, Y => n103);
   U125 : INVX2 port map( A => n81, Y => n106);
   U127 : INVX2 port map( A => n82, Y => n113);
   U131 : INVX2 port map( A => n78, Y => n118);
   U135 : INVX2 port map( A => n54, Y => n121);
   U137 : INVX2 port map( A => n171, Y => n125);
   U138 : INVX2 port map( A => n101, Y => n131);
   U144 : INVX2 port map( A => n102, Y => n136);
   U151 : INVX2 port map( A => n97, Y => n139);
   U158 : INVX2 port map( A => n98, Y => n145);
   U161 : INVX2 port map( A => n94, Y => n148);
   U165 : INVX2 port map( A => n87, Y => n152);
   U168 : INVX2 port map( A => n88, Y => n153);
   U170 : INVX2 port map( A => n150, Y => n164);
   U179 : INVX2 port map( A => n3, Y => n168);
   U180 : INVX2 port map( A => n1, Y => n175);
   U181 : INVX2 port map( A => n119, Y => n181);
   U182 : INVX2 port map( A => n68, Y => n188);
   U183 : INVX2 port map( A => n172, Y => n191);
   U185 : INVX2 port map( A => n48, Y => n192);
   U186 : INVX2 port map( A => n149, Y => n211);
   U188 : INVX2 port map( A => n274, Y => n213);
   U191 : INVX2 port map( A => n141, Y => init_math);
   U195 : INVX2 port map( A => n49, Y => n215);
   U196 : INVX2 port map( A => n69, Y => n216);
   U198 : INVX2 port map( A => counter_4_port, Y => n217);
   U202 : INVX2 port map( A => n176, Y => n218);
   U203 : INVX2 port map( A => n127, Y => n219);
   U206 : INVX2 port map( A => state_2_port, Y => n220);
   U208 : INVX2 port map( A => state_0_port, Y => n221);
   U211 : INVX2 port map( A => state_1_port, Y => n222);
   U213 : INVX2 port map( A => opp_0_port, Y => n223);
   U220 : INVX2 port map( A => opp_1_port, Y => n224);
   U228 : INVX2 port map( A => n165, Y => n225);
   U234 : INVX2 port map( A => opp_6_port, Y => n226);
   U238 : INVX2 port map( A => opp_7_port, Y => n227);
   U241 : INVX2 port map( A => n169, Y => n228);
   U243 : INVX2 port map( A => opp_13_port, Y => n275);
   U244 : INVX2 port map( A => opp_14_port, Y => n292);
   U246 : INVX2 port map( A => counter_3_port, Y => n299_port);
   U248 : INVX2 port map( A => counter_0_port, Y => n301_port);
   U265 : INVX2 port map( A => counter_1_port, Y => n302_port);
   U270 : INVX2 port map( A => counter_2_port, Y => n303_port);
   U272 : INVX2 port map( A => addr_0_port, Y => n304_port);
   U273 : INVX2 port map( A => addr_1_port, Y => n305_port);
   U275 : INVX2 port map( A => addr_2_port, Y => n306_port);
   U279 : INVX2 port map( A => addr_3_port, Y => n307_port);
   U280 : INVX2 port map( A => addr_4_port, Y => n308_port);
   U281 : INVX2 port map( A => addr_5_port, Y => n309_port);
   U282 : INVX2 port map( A => addr_6_port, Y => n310_port);
   U283 : INVX2 port map( A => addr_7_port, Y => n311_port);
   U284 : INVX2 port map( A => addr_8_port, Y => n313);
   U285 : INVX2 port map( A => addr_9_port, Y => n315_port);
   U286 : INVX2 port map( A => addr_10_port, Y => n316_port);
   U287 : INVX2 port map( A => addr_11_port, Y => n317_port);
   U288 : INVX2 port map( A => addr_12_port, Y => n318);
   U289 : INVX2 port map( A => addr_13_port, Y => n319);
   U290 : INVX2 port map( A => addr_14_port, Y => n320);
   U291 : INVX2 port map( A => re, Y => n321);
   U292 : INVX2 port map( A => rast_strb, Y => n322);
   U293 : INVX2 port map( A => rast_index(2), Y => n323);
   U294 : INVX2 port map( A => rast_index(3), Y => n325);
   U340 : INVX2 port map( A => rast_index(0), Y => n327);
   U341 : INVX2 port map( A => math_done, Y => n332);

end SYN_struct;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity coordinate_buffer is

   port( strb_cor : in std_logic;  databus_out : in std_logic_vector (15 downto
         0);  clk, sel : in std_logic;  point : out std_logic_vector (47 downto
         0));

end coordinate_buffer;

architecture SYN_behavorial of coordinate_buffer is

   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal regg_95_port, regg_94_port, regg_93_port, regg_92_port, regg_91_port,
      regg_90_port, regg_89_port, regg_88_port, regg_87_port, regg_86_port, 
      regg_85_port, regg_84_port, regg_83_port, regg_82_port, regg_81_port, 
      regg_80_port, regg_79_port, regg_78_port, regg_77_port, regg_76_port, 
      regg_75_port, regg_74_port, regg_73_port, regg_72_port, regg_71_port, 
      regg_70_port, regg_69_port, regg_68_port, regg_67_port, regg_66_port, 
      regg_65_port, regg_64_port, regg_63_port, regg_62_port, regg_61_port, 
      regg_60_port, regg_59_port, regg_58_port, regg_57_port, regg_56_port, 
      regg_55_port, regg_54_port, regg_53_port, regg_52_port, regg_51_port, 
      regg_50_port, regg_49_port, regg_48_port, regg_47_port, regg_46_port, 
      regg_45_port, regg_44_port, regg_43_port, regg_42_port, regg_41_port, 
      regg_40_port, regg_39_port, regg_38_port, regg_37_port, regg_36_port, 
      regg_35_port, regg_34_port, regg_33_port, regg_32_port, regg_31_port, 
      regg_30_port, regg_29_port, regg_28_port, regg_27_port, regg_26_port, 
      regg_25_port, regg_24_port, regg_23_port, regg_22_port, regg_21_port, 
      regg_20_port, regg_19_port, regg_18_port, regg_17_port, regg_16_port, 
      regg_15_port, regg_14_port, regg_13_port, regg_12_port, regg_11_port, 
      regg_10_port, regg_9_port, regg_8_port, regg_7_port, regg_6_port, 
      regg_5_port, regg_4_port, regg_3_port, regg_2_port, regg_1_port, 
      regg_0_port, n8, n15, n22, n29, n36, n43, n50, n57, n64, n71, n78, n85, 
      n92, n99, n106, n113, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, 
      n13, n14, n16, n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n30
      , n31, n32, n33, n34, n35, n37, n38, n39, n40, n41, n42, n44, n45, n46, 
      n47, n48, n49, n51, n52, n53, n54, n55, n56, n58, n59, n60, n61, n62, n63
      , n65, n66, n67, n68, n69, n70, n72, n73, n74, n75, n76, n77, n79, n80, 
      n81, n82, n83, n84, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97
      , n98, n100, n101, n102, n103, n104, n105, n107, n108, n109, n110, n111, 
      n112, n114, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244 : 
      std_logic;

begin
   
   regg_reg_15_inst : DFFPOSX1 port map( D => n210, CLK => clk, Q => 
                           regg_15_port);
   regg_reg_31_inst : DFFPOSX1 port map( D => n209, CLK => clk, Q => 
                           regg_31_port);
   regg_reg_47_inst : DFFPOSX1 port map( D => n208, CLK => clk, Q => 
                           regg_47_port);
   regg_reg_63_inst : DFFPOSX1 port map( D => n207, CLK => clk, Q => 
                           regg_63_port);
   regg_reg_79_inst : DFFPOSX1 port map( D => n206, CLK => clk, Q => 
                           regg_79_port);
   regg_reg_95_inst : DFFPOSX1 port map( D => n205, CLK => clk, Q => 
                           regg_95_port);
   regg_reg_14_inst : DFFPOSX1 port map( D => n204, CLK => clk, Q => 
                           regg_14_port);
   regg_reg_30_inst : DFFPOSX1 port map( D => n203, CLK => clk, Q => 
                           regg_30_port);
   regg_reg_46_inst : DFFPOSX1 port map( D => n202, CLK => clk, Q => 
                           regg_46_port);
   regg_reg_62_inst : DFFPOSX1 port map( D => n201, CLK => clk, Q => 
                           regg_62_port);
   regg_reg_78_inst : DFFPOSX1 port map( D => n200, CLK => clk, Q => 
                           regg_78_port);
   regg_reg_94_inst : DFFPOSX1 port map( D => n199, CLK => clk, Q => 
                           regg_94_port);
   regg_reg_13_inst : DFFPOSX1 port map( D => n198, CLK => clk, Q => 
                           regg_13_port);
   regg_reg_29_inst : DFFPOSX1 port map( D => n197, CLK => clk, Q => 
                           regg_29_port);
   regg_reg_45_inst : DFFPOSX1 port map( D => n196, CLK => clk, Q => 
                           regg_45_port);
   regg_reg_61_inst : DFFPOSX1 port map( D => n195, CLK => clk, Q => 
                           regg_61_port);
   regg_reg_77_inst : DFFPOSX1 port map( D => n194, CLK => clk, Q => 
                           regg_77_port);
   regg_reg_93_inst : DFFPOSX1 port map( D => n193, CLK => clk, Q => 
                           regg_93_port);
   regg_reg_12_inst : DFFPOSX1 port map( D => n192, CLK => clk, Q => 
                           regg_12_port);
   regg_reg_28_inst : DFFPOSX1 port map( D => n191, CLK => clk, Q => 
                           regg_28_port);
   regg_reg_44_inst : DFFPOSX1 port map( D => n190, CLK => clk, Q => 
                           regg_44_port);
   regg_reg_60_inst : DFFPOSX1 port map( D => n189, CLK => clk, Q => 
                           regg_60_port);
   regg_reg_76_inst : DFFPOSX1 port map( D => n188, CLK => clk, Q => 
                           regg_76_port);
   regg_reg_92_inst : DFFPOSX1 port map( D => n187, CLK => clk, Q => 
                           regg_92_port);
   regg_reg_11_inst : DFFPOSX1 port map( D => n186, CLK => clk, Q => 
                           regg_11_port);
   regg_reg_27_inst : DFFPOSX1 port map( D => n185, CLK => clk, Q => 
                           regg_27_port);
   regg_reg_43_inst : DFFPOSX1 port map( D => n184, CLK => clk, Q => 
                           regg_43_port);
   regg_reg_59_inst : DFFPOSX1 port map( D => n183, CLK => clk, Q => 
                           regg_59_port);
   regg_reg_75_inst : DFFPOSX1 port map( D => n182, CLK => clk, Q => 
                           regg_75_port);
   regg_reg_91_inst : DFFPOSX1 port map( D => n181, CLK => clk, Q => 
                           regg_91_port);
   regg_reg_10_inst : DFFPOSX1 port map( D => n180, CLK => clk, Q => 
                           regg_10_port);
   regg_reg_26_inst : DFFPOSX1 port map( D => n179, CLK => clk, Q => 
                           regg_26_port);
   regg_reg_42_inst : DFFPOSX1 port map( D => n178, CLK => clk, Q => 
                           regg_42_port);
   regg_reg_58_inst : DFFPOSX1 port map( D => n177, CLK => clk, Q => 
                           regg_58_port);
   regg_reg_74_inst : DFFPOSX1 port map( D => n176, CLK => clk, Q => 
                           regg_74_port);
   regg_reg_90_inst : DFFPOSX1 port map( D => n175, CLK => clk, Q => 
                           regg_90_port);
   regg_reg_9_inst : DFFPOSX1 port map( D => n174, CLK => clk, Q => regg_9_port
                           );
   regg_reg_25_inst : DFFPOSX1 port map( D => n173, CLK => clk, Q => 
                           regg_25_port);
   regg_reg_41_inst : DFFPOSX1 port map( D => n172, CLK => clk, Q => 
                           regg_41_port);
   regg_reg_57_inst : DFFPOSX1 port map( D => n171, CLK => clk, Q => 
                           regg_57_port);
   regg_reg_73_inst : DFFPOSX1 port map( D => n170, CLK => clk, Q => 
                           regg_73_port);
   regg_reg_89_inst : DFFPOSX1 port map( D => n169, CLK => clk, Q => 
                           regg_89_port);
   regg_reg_8_inst : DFFPOSX1 port map( D => n168, CLK => clk, Q => regg_8_port
                           );
   regg_reg_24_inst : DFFPOSX1 port map( D => n167, CLK => clk, Q => 
                           regg_24_port);
   regg_reg_40_inst : DFFPOSX1 port map( D => n166, CLK => clk, Q => 
                           regg_40_port);
   regg_reg_56_inst : DFFPOSX1 port map( D => n165, CLK => clk, Q => 
                           regg_56_port);
   regg_reg_72_inst : DFFPOSX1 port map( D => n164, CLK => clk, Q => 
                           regg_72_port);
   regg_reg_88_inst : DFFPOSX1 port map( D => n163, CLK => clk, Q => 
                           regg_88_port);
   regg_reg_7_inst : DFFPOSX1 port map( D => n162, CLK => clk, Q => regg_7_port
                           );
   regg_reg_23_inst : DFFPOSX1 port map( D => n161, CLK => clk, Q => 
                           regg_23_port);
   regg_reg_39_inst : DFFPOSX1 port map( D => n160, CLK => clk, Q => 
                           regg_39_port);
   regg_reg_55_inst : DFFPOSX1 port map( D => n159, CLK => clk, Q => 
                           regg_55_port);
   regg_reg_71_inst : DFFPOSX1 port map( D => n158, CLK => clk, Q => 
                           regg_71_port);
   regg_reg_87_inst : DFFPOSX1 port map( D => n157, CLK => clk, Q => 
                           regg_87_port);
   regg_reg_6_inst : DFFPOSX1 port map( D => n156, CLK => clk, Q => regg_6_port
                           );
   regg_reg_22_inst : DFFPOSX1 port map( D => n155, CLK => clk, Q => 
                           regg_22_port);
   regg_reg_38_inst : DFFPOSX1 port map( D => n154, CLK => clk, Q => 
                           regg_38_port);
   regg_reg_54_inst : DFFPOSX1 port map( D => n153, CLK => clk, Q => 
                           regg_54_port);
   regg_reg_70_inst : DFFPOSX1 port map( D => n152, CLK => clk, Q => 
                           regg_70_port);
   regg_reg_86_inst : DFFPOSX1 port map( D => n151, CLK => clk, Q => 
                           regg_86_port);
   regg_reg_5_inst : DFFPOSX1 port map( D => n150, CLK => clk, Q => regg_5_port
                           );
   regg_reg_21_inst : DFFPOSX1 port map( D => n149, CLK => clk, Q => 
                           regg_21_port);
   regg_reg_37_inst : DFFPOSX1 port map( D => n148, CLK => clk, Q => 
                           regg_37_port);
   regg_reg_53_inst : DFFPOSX1 port map( D => n147, CLK => clk, Q => 
                           regg_53_port);
   regg_reg_69_inst : DFFPOSX1 port map( D => n146, CLK => clk, Q => 
                           regg_69_port);
   regg_reg_85_inst : DFFPOSX1 port map( D => n145, CLK => clk, Q => 
                           regg_85_port);
   regg_reg_4_inst : DFFPOSX1 port map( D => n144, CLK => clk, Q => regg_4_port
                           );
   regg_reg_20_inst : DFFPOSX1 port map( D => n143, CLK => clk, Q => 
                           regg_20_port);
   regg_reg_36_inst : DFFPOSX1 port map( D => n142, CLK => clk, Q => 
                           regg_36_port);
   regg_reg_52_inst : DFFPOSX1 port map( D => n141, CLK => clk, Q => 
                           regg_52_port);
   regg_reg_68_inst : DFFPOSX1 port map( D => n140, CLK => clk, Q => 
                           regg_68_port);
   regg_reg_84_inst : DFFPOSX1 port map( D => n139, CLK => clk, Q => 
                           regg_84_port);
   regg_reg_3_inst : DFFPOSX1 port map( D => n138, CLK => clk, Q => regg_3_port
                           );
   regg_reg_19_inst : DFFPOSX1 port map( D => n137, CLK => clk, Q => 
                           regg_19_port);
   regg_reg_35_inst : DFFPOSX1 port map( D => n136, CLK => clk, Q => 
                           regg_35_port);
   regg_reg_51_inst : DFFPOSX1 port map( D => n135, CLK => clk, Q => 
                           regg_51_port);
   regg_reg_67_inst : DFFPOSX1 port map( D => n134, CLK => clk, Q => 
                           regg_67_port);
   regg_reg_83_inst : DFFPOSX1 port map( D => n133, CLK => clk, Q => 
                           regg_83_port);
   regg_reg_2_inst : DFFPOSX1 port map( D => n132, CLK => clk, Q => regg_2_port
                           );
   regg_reg_18_inst : DFFPOSX1 port map( D => n131, CLK => clk, Q => 
                           regg_18_port);
   regg_reg_34_inst : DFFPOSX1 port map( D => n130, CLK => clk, Q => 
                           regg_34_port);
   regg_reg_50_inst : DFFPOSX1 port map( D => n129, CLK => clk, Q => 
                           regg_50_port);
   regg_reg_66_inst : DFFPOSX1 port map( D => n128, CLK => clk, Q => 
                           regg_66_port);
   regg_reg_82_inst : DFFPOSX1 port map( D => n127, CLK => clk, Q => 
                           regg_82_port);
   regg_reg_1_inst : DFFPOSX1 port map( D => n126, CLK => clk, Q => regg_1_port
                           );
   regg_reg_17_inst : DFFPOSX1 port map( D => n125, CLK => clk, Q => 
                           regg_17_port);
   regg_reg_33_inst : DFFPOSX1 port map( D => n124, CLK => clk, Q => 
                           regg_33_port);
   regg_reg_49_inst : DFFPOSX1 port map( D => n123, CLK => clk, Q => 
                           regg_49_port);
   regg_reg_65_inst : DFFPOSX1 port map( D => n122, CLK => clk, Q => 
                           regg_65_port);
   regg_reg_81_inst : DFFPOSX1 port map( D => n121, CLK => clk, Q => 
                           regg_81_port);
   regg_reg_0_inst : DFFPOSX1 port map( D => n120, CLK => clk, Q => regg_0_port
                           );
   regg_reg_16_inst : DFFPOSX1 port map( D => n119, CLK => clk, Q => 
                           regg_16_port);
   regg_reg_32_inst : DFFPOSX1 port map( D => n118, CLK => clk, Q => 
                           regg_32_port);
   regg_reg_48_inst : DFFPOSX1 port map( D => n117, CLK => clk, Q => 
                           regg_48_port);
   regg_reg_64_inst : DFFPOSX1 port map( D => n116, CLK => clk, Q => 
                           regg_64_port);
   regg_reg_80_inst : DFFPOSX1 port map( D => n115, CLK => clk, Q => 
                           regg_80_port);
   U8 : NAND2X1 port map( A => databus_out(0), B => n11, Y => n8);
   U15 : NAND2X1 port map( A => databus_out(1), B => n13, Y => n15);
   U22 : NAND2X1 port map( A => databus_out(2), B => n10, Y => n22);
   U29 : NAND2X1 port map( A => databus_out(3), B => n12, Y => n29);
   U36 : NAND2X1 port map( A => databus_out(4), B => n14, Y => n36);
   U43 : NAND2X1 port map( A => databus_out(5), B => n11, Y => n43);
   U50 : NAND2X1 port map( A => databus_out(6), B => n13, Y => n50);
   U57 : NAND2X1 port map( A => databus_out(7), B => n11, Y => n57);
   U64 : NAND2X1 port map( A => databus_out(8), B => n16, Y => n64);
   U71 : NAND2X1 port map( A => databus_out(9), B => n13, Y => n71);
   U78 : NAND2X1 port map( A => databus_out(10), B => n9, Y => n78);
   U85 : NAND2X1 port map( A => databus_out(11), B => n9, Y => n85);
   U92 : NAND2X1 port map( A => databus_out(12), B => n9, Y => n92);
   U99 : NAND2X1 port map( A => databus_out(13), B => n10, Y => n99);
   U106 : NAND2X1 port map( A => databus_out(14), B => n12, Y => n106);
   U114 : NAND2X1 port map( A => databus_out(15), B => n9, Y => n113);
   U2 : INVX2 port map( A => n4, Y => n2);
   U3 : INVX1 port map( A => n40, Y => n1);
   U4 : BUFX4 port map( A => sel, Y => n3);
   U5 : INVX2 port map( A => sel, Y => n40);
   U6 : MUX2X1 port map( B => n111, A => n108, S => n40, Y => point(9));
   U7 : MUX2X1 port map( B => n237, A => n234, S => n40, Y => point(30));
   U9 : MUX2X1 port map( B => n232, A => n229, S => n40, Y => point(13));
   U10 : MUX2X1 port map( B => n213, A => n114, S => n40, Y => point(26));
   U11 : BUFX4 port map( A => sel, Y => n4);
   U12 : MUX2X1 port map( B => n62, A => n59, S => n2, Y => point(2));
   U13 : INVX2 port map( A => n25, Y => n10);
   U14 : INVX2 port map( A => n19, Y => n16);
   U16 : INVX2 port map( A => n20, Y => n14);
   U17 : INVX2 port map( A => n21, Y => n13);
   U18 : INVX2 port map( A => n24, Y => n11);
   U19 : INVX2 port map( A => n23, Y => n12);
   U20 : INVX2 port map( A => n26, Y => n9);
   U21 : BUFX2 port map( A => n37, Y => n19);
   U23 : BUFX2 port map( A => n37, Y => n20);
   U24 : BUFX2 port map( A => n37, Y => n21);
   U25 : BUFX2 port map( A => n37, Y => n23);
   U26 : BUFX2 port map( A => n37, Y => n24);
   U27 : BUFX2 port map( A => n37, Y => n25);
   U28 : BUFX2 port map( A => n37, Y => n26);
   U30 : BUFX2 port map( A => n37, Y => n17);
   U31 : BUFX2 port map( A => n37, Y => n18);
   U32 : BUFX2 port map( A => n17, Y => n27);
   U33 : BUFX2 port map( A => n17, Y => n28);
   U34 : BUFX2 port map( A => n17, Y => n30);
   U35 : BUFX2 port map( A => n37, Y => n31);
   U37 : BUFX2 port map( A => n37, Y => n32);
   U38 : BUFX2 port map( A => n37, Y => n33);
   U39 : BUFX2 port map( A => n37, Y => n34);
   U40 : BUFX2 port map( A => n37, Y => n35);
   U41 : INVX2 port map( A => strb_cor, Y => n37);
   U42 : INVX4 port map( A => n6, Y => point(31));
   U44 : INVX4 port map( A => n7, Y => point(15));
   U45 : INVX4 port map( A => n5, Y => point(47));
   U46 : MUX2X1 port map( B => regg_95_port, A => regg_47_port, S => n38, Y => 
                           n5);
   U47 : INVX1 port map( A => regg_95_port, Y => n239);
   U48 : INVX1 port map( A => regg_47_port, Y => n242);
   U49 : INVX4 port map( A => sel, Y => n41);
   U51 : MUX2X1 port map( B => regg_31_port, A => regg_79_port, S => n2, Y => 
                           n6);
   U52 : INVX1 port map( A => regg_31_port, Y => n243);
   U53 : INVX1 port map( A => regg_79_port, Y => n240);
   U54 : MUX2X1 port map( B => regg_15_port, A => regg_63_port, S => n40, Y => 
                           n7);
   U55 : INVX1 port map( A => regg_15_port, Y => n244);
   U56 : INVX1 port map( A => regg_63_port, Y => n241);
   U58 : INVX8 port map( A => n41, Y => n38);
   U59 : INVX8 port map( A => n41, Y => n39);
   U60 : INVX2 port map( A => regg_48_port, Y => n45);
   U61 : INVX2 port map( A => regg_0_port, Y => n48);
   U62 : MUX2X1 port map( B => n45, A => n48, S => n38, Y => point(0));
   U63 : INVX2 port map( A => regg_49_port, Y => n52);
   U65 : INVX2 port map( A => regg_1_port, Y => n55);
   U66 : MUX2X1 port map( B => n52, A => n55, S => n38, Y => point(1));
   U67 : INVX2 port map( A => regg_50_port, Y => n59);
   U68 : INVX2 port map( A => regg_2_port, Y => n62);
   U69 : INVX2 port map( A => regg_51_port, Y => n66);
   U70 : INVX2 port map( A => regg_3_port, Y => n69);
   U72 : MUX2X1 port map( B => n66, A => n69, S => n38, Y => point(3));
   U73 : INVX2 port map( A => regg_52_port, Y => n73);
   U74 : INVX2 port map( A => regg_4_port, Y => n76);
   U75 : MUX2X1 port map( B => n73, A => n76, S => n38, Y => point(4));
   U76 : INVX2 port map( A => regg_53_port, Y => n80);
   U77 : INVX2 port map( A => regg_5_port, Y => n83);
   U79 : MUX2X1 port map( B => n80, A => n83, S => n38, Y => point(5));
   U80 : INVX2 port map( A => regg_54_port, Y => n87);
   U81 : INVX2 port map( A => regg_6_port, Y => n90);
   U82 : MUX2X1 port map( B => n87, A => n90, S => n38, Y => point(6));
   U83 : INVX2 port map( A => regg_55_port, Y => n94);
   U84 : INVX2 port map( A => regg_7_port, Y => n97);
   U86 : MUX2X1 port map( B => n94, A => n97, S => n38, Y => point(7));
   U87 : INVX2 port map( A => regg_56_port, Y => n101);
   U88 : INVX2 port map( A => regg_8_port, Y => n104);
   U89 : MUX2X1 port map( B => n101, A => n104, S => n39, Y => point(8));
   U90 : INVX2 port map( A => regg_57_port, Y => n108);
   U91 : INVX2 port map( A => regg_9_port, Y => n111);
   U93 : INVX2 port map( A => regg_58_port, Y => n211);
   U94 : INVX2 port map( A => regg_10_port, Y => n214);
   U95 : MUX2X1 port map( B => n211, A => n214, S => n38, Y => point(10));
   U96 : INVX2 port map( A => regg_59_port, Y => n217);
   U97 : INVX2 port map( A => regg_11_port, Y => n220);
   U98 : MUX2X1 port map( B => n217, A => n220, S => n4, Y => point(11));
   U100 : INVX2 port map( A => regg_60_port, Y => n223);
   U101 : INVX2 port map( A => regg_12_port, Y => n226);
   U102 : MUX2X1 port map( B => n223, A => n226, S => n3, Y => point(12));
   U103 : INVX2 port map( A => regg_61_port, Y => n229);
   U104 : INVX2 port map( A => regg_13_port, Y => n232);
   U105 : INVX2 port map( A => regg_62_port, Y => n235);
   U107 : INVX2 port map( A => regg_14_port, Y => n238);
   U108 : MUX2X1 port map( B => n235, A => n238, S => n39, Y => point(14));
   U109 : INVX2 port map( A => regg_64_port, Y => n44);
   U110 : INVX2 port map( A => regg_16_port, Y => n47);
   U111 : MUX2X1 port map( B => n44, A => n47, S => n38, Y => point(16));
   U112 : INVX2 port map( A => regg_65_port, Y => n51);
   U113 : INVX2 port map( A => regg_17_port, Y => n54);
   U115 : MUX2X1 port map( B => n51, A => n54, S => n38, Y => point(17));
   U116 : INVX2 port map( A => regg_66_port, Y => n58);
   U117 : INVX2 port map( A => regg_18_port, Y => n61);
   U118 : MUX2X1 port map( B => n58, A => n61, S => n38, Y => point(18));
   U119 : INVX2 port map( A => regg_67_port, Y => n65);
   U120 : INVX2 port map( A => regg_19_port, Y => n68);
   U121 : MUX2X1 port map( B => n65, A => n68, S => n38, Y => point(19));
   U122 : INVX2 port map( A => regg_68_port, Y => n72);
   U123 : INVX2 port map( A => regg_20_port, Y => n75);
   U124 : MUX2X1 port map( B => n72, A => n75, S => n39, Y => point(20));
   U125 : INVX2 port map( A => regg_69_port, Y => n79);
   U126 : INVX2 port map( A => regg_21_port, Y => n82);
   U127 : MUX2X1 port map( B => n79, A => n82, S => n39, Y => point(21));
   U128 : INVX2 port map( A => regg_70_port, Y => n86);
   U129 : INVX2 port map( A => regg_22_port, Y => n89);
   U130 : MUX2X1 port map( B => n86, A => n89, S => n39, Y => point(22));
   U131 : INVX2 port map( A => regg_71_port, Y => n93);
   U132 : INVX2 port map( A => regg_23_port, Y => n96);
   U133 : MUX2X1 port map( B => n93, A => n96, S => n38, Y => point(23));
   U134 : INVX2 port map( A => regg_72_port, Y => n100);
   U135 : INVX2 port map( A => regg_24_port, Y => n103);
   U136 : MUX2X1 port map( B => n100, A => n103, S => n3, Y => point(24));
   U137 : INVX2 port map( A => regg_73_port, Y => n107);
   U138 : INVX2 port map( A => regg_25_port, Y => n110);
   U139 : MUX2X1 port map( B => n107, A => n110, S => n4, Y => point(25));
   U140 : INVX2 port map( A => regg_74_port, Y => n114);
   U141 : INVX2 port map( A => regg_26_port, Y => n213);
   U142 : INVX2 port map( A => regg_75_port, Y => n216);
   U143 : INVX2 port map( A => regg_27_port, Y => n219);
   U144 : MUX2X1 port map( B => n216, A => n219, S => n39, Y => point(27));
   U145 : INVX2 port map( A => regg_76_port, Y => n222);
   U146 : INVX2 port map( A => regg_28_port, Y => n225);
   U147 : MUX2X1 port map( B => n222, A => n225, S => n4, Y => point(28));
   U148 : INVX2 port map( A => regg_77_port, Y => n228);
   U149 : INVX2 port map( A => regg_29_port, Y => n231);
   U150 : MUX2X1 port map( B => n228, A => n231, S => n39, Y => point(29));
   U151 : INVX2 port map( A => regg_78_port, Y => n234);
   U152 : INVX2 port map( A => regg_30_port, Y => n237);
   U153 : INVX2 port map( A => regg_80_port, Y => n42);
   U154 : INVX2 port map( A => regg_32_port, Y => n46);
   U155 : MUX2X1 port map( B => n42, A => n46, S => n38, Y => point(32));
   U156 : INVX2 port map( A => regg_81_port, Y => n49);
   U157 : INVX2 port map( A => regg_33_port, Y => n53);
   U158 : MUX2X1 port map( B => n49, A => n53, S => n38, Y => point(33));
   U159 : INVX2 port map( A => regg_82_port, Y => n56);
   U160 : INVX2 port map( A => regg_34_port, Y => n60);
   U161 : MUX2X1 port map( B => n56, A => n60, S => n38, Y => point(34));
   U162 : INVX2 port map( A => regg_83_port, Y => n63);
   U163 : INVX2 port map( A => regg_35_port, Y => n67);
   U164 : MUX2X1 port map( B => n63, A => n67, S => n38, Y => point(35));
   U165 : INVX2 port map( A => regg_84_port, Y => n70);
   U166 : INVX2 port map( A => regg_36_port, Y => n74);
   U167 : MUX2X1 port map( B => n70, A => n74, S => n39, Y => point(36));
   U168 : INVX2 port map( A => regg_85_port, Y => n77);
   U169 : INVX2 port map( A => regg_37_port, Y => n81);
   U170 : MUX2X1 port map( B => n77, A => n81, S => n38, Y => point(37));
   U171 : INVX2 port map( A => regg_86_port, Y => n84);
   U172 : INVX2 port map( A => regg_38_port, Y => n88);
   U173 : MUX2X1 port map( B => n84, A => n88, S => n3, Y => point(38));
   U174 : INVX2 port map( A => regg_87_port, Y => n91);
   U175 : INVX2 port map( A => regg_39_port, Y => n95);
   U176 : MUX2X1 port map( B => n91, A => n95, S => n3, Y => point(39));
   U177 : INVX2 port map( A => regg_88_port, Y => n98);
   U178 : INVX2 port map( A => regg_40_port, Y => n102);
   U179 : MUX2X1 port map( B => n98, A => n102, S => n3, Y => point(40));
   U180 : INVX2 port map( A => regg_89_port, Y => n105);
   U181 : INVX2 port map( A => regg_41_port, Y => n109);
   U182 : MUX2X1 port map( B => n105, A => n109, S => n3, Y => point(41));
   U183 : INVX2 port map( A => regg_90_port, Y => n112);
   U184 : INVX2 port map( A => regg_42_port, Y => n212);
   U185 : MUX2X1 port map( B => n112, A => n212, S => n39, Y => point(42));
   U186 : INVX2 port map( A => regg_91_port, Y => n215);
   U187 : INVX2 port map( A => regg_43_port, Y => n218);
   U188 : MUX2X1 port map( B => n215, A => n218, S => n4, Y => point(43));
   U189 : INVX2 port map( A => regg_92_port, Y => n221);
   U190 : INVX2 port map( A => regg_44_port, Y => n224);
   U191 : MUX2X1 port map( B => n221, A => n224, S => n1, Y => point(44));
   U192 : INVX2 port map( A => regg_93_port, Y => n227);
   U193 : INVX2 port map( A => regg_45_port, Y => n230);
   U194 : MUX2X1 port map( B => n227, A => n230, S => n39, Y => point(45));
   U195 : INVX2 port map( A => regg_94_port, Y => n233);
   U196 : INVX2 port map( A => regg_46_port, Y => n236);
   U197 : MUX2X1 port map( B => n233, A => n236, S => n38, Y => point(46));
   U198 : OAI22X1 port map( A => n42, B => n13, C => n17, D => n44, Y => n115);
   U199 : OAI22X1 port map( A => n44, B => n12, C => n17, D => n45, Y => n116);
   U200 : OAI22X1 port map( A => n45, B => n10, C => n17, D => n46, Y => n117);
   U201 : OAI22X1 port map( A => n46, B => n13, C => n18, D => n47, Y => n118);
   U202 : OAI22X1 port map( A => n47, B => n11, C => n18, D => n48, Y => n119);
   U203 : OAI21X1 port map( A => n48, B => n9, C => n8, Y => n120);
   U204 : OAI22X1 port map( A => n49, B => n16, C => n18, D => n51, Y => n121);
   U205 : OAI22X1 port map( A => n51, B => n14, C => n19, D => n52, Y => n122);
   U206 : OAI22X1 port map( A => n52, B => n16, C => n19, D => n53, Y => n123);
   U207 : OAI22X1 port map( A => n53, B => n16, C => n19, D => n54, Y => n124);
   U208 : OAI22X1 port map( A => n54, B => n16, C => n20, D => n55, Y => n125);
   U209 : OAI21X1 port map( A => n55, B => n9, C => n15, Y => n126);
   U210 : OAI22X1 port map( A => n56, B => n16, C => n20, D => n58, Y => n127);
   U211 : OAI22X1 port map( A => n58, B => n16, C => n20, D => n59, Y => n128);
   U212 : OAI22X1 port map( A => n59, B => n16, C => n21, D => n60, Y => n129);
   U213 : OAI22X1 port map( A => n60, B => n16, C => n21, D => n61, Y => n130);
   U214 : OAI22X1 port map( A => n61, B => n16, C => n21, D => n62, Y => n131);
   U215 : OAI21X1 port map( A => n62, B => n9, C => n22, Y => n132);
   U216 : OAI22X1 port map( A => n63, B => n16, C => n23, D => n65, Y => n133);
   U217 : OAI22X1 port map( A => n65, B => n16, C => n23, D => n66, Y => n134);
   U218 : OAI22X1 port map( A => n66, B => n16, C => n23, D => n67, Y => n135);
   U219 : OAI22X1 port map( A => n67, B => n16, C => n24, D => n68, Y => n136);
   U220 : OAI22X1 port map( A => n68, B => n16, C => n24, D => n69, Y => n137);
   U221 : OAI21X1 port map( A => n69, B => n9, C => n29, Y => n138);
   U222 : OAI22X1 port map( A => n70, B => n14, C => n24, D => n72, Y => n139);
   U223 : OAI22X1 port map( A => n72, B => n14, C => n25, D => n73, Y => n140);
   U224 : OAI22X1 port map( A => n73, B => n14, C => n25, D => n74, Y => n141);
   U225 : OAI22X1 port map( A => n74, B => n14, C => n25, D => n75, Y => n142);
   U226 : OAI22X1 port map( A => n75, B => n14, C => n26, D => n76, Y => n143);
   U227 : OAI21X1 port map( A => n76, B => n10, C => n36, Y => n144);
   U228 : OAI22X1 port map( A => n77, B => n14, C => n26, D => n79, Y => n145);
   U229 : OAI22X1 port map( A => n79, B => n14, C => n26, D => n80, Y => n146);
   U230 : OAI22X1 port map( A => n80, B => n14, C => n27, D => n81, Y => n147);
   U231 : OAI22X1 port map( A => n81, B => n14, C => n27, D => n82, Y => n148);
   U232 : OAI22X1 port map( A => n82, B => n14, C => n27, D => n83, Y => n149);
   U233 : OAI21X1 port map( A => n83, B => n9, C => n43, Y => n150);
   U234 : OAI22X1 port map( A => n84, B => n14, C => n27, D => n86, Y => n151);
   U235 : OAI22X1 port map( A => n86, B => n14, C => n27, D => n87, Y => n152);
   U236 : OAI22X1 port map( A => n87, B => n14, C => n27, D => n88, Y => n153);
   U237 : OAI22X1 port map( A => n88, B => n13, C => n27, D => n89, Y => n154);
   U238 : OAI22X1 port map( A => n89, B => n13, C => n28, D => n90, Y => n155);
   U239 : OAI21X1 port map( A => n90, B => n9, C => n50, Y => n156);
   U240 : OAI22X1 port map( A => n91, B => n13, C => n28, D => n93, Y => n157);
   U241 : OAI22X1 port map( A => n93, B => n13, C => n28, D => n94, Y => n158);
   U242 : OAI22X1 port map( A => n94, B => n13, C => n28, D => n95, Y => n159);
   U243 : OAI22X1 port map( A => n95, B => n13, C => n28, D => n96, Y => n160);
   U244 : OAI22X1 port map( A => n96, B => n13, C => n28, D => n97, Y => n161);
   U245 : OAI21X1 port map( A => n97, B => n9, C => n57, Y => n162);
   U246 : OAI22X1 port map( A => n98, B => n13, C => n28, D => n100, Y => n163)
                           ;
   U247 : OAI22X1 port map( A => n100, B => n13, C => n30, D => n101, Y => n164
                           );
   U248 : OAI22X1 port map( A => n101, B => n13, C => n30, D => n102, Y => n165
                           );
   U249 : OAI22X1 port map( A => n102, B => n13, C => n30, D => n103, Y => n166
                           );
   U250 : OAI22X1 port map( A => n103, B => n13, C => n30, D => n104, Y => n167
                           );
   U251 : OAI21X1 port map( A => n104, B => n10, C => n64, Y => n168);
   U252 : OAI22X1 port map( A => n105, B => n12, C => n30, D => n107, Y => n169
                           );
   U253 : OAI22X1 port map( A => n107, B => n12, C => n30, D => n108, Y => n170
                           );
   U254 : OAI22X1 port map( A => n108, B => n12, C => n30, D => n109, Y => n171
                           );
   U255 : OAI22X1 port map( A => n109, B => n12, C => n31, D => n110, Y => n172
                           );
   U256 : OAI22X1 port map( A => n110, B => n12, C => n31, D => n111, Y => n173
                           );
   U257 : OAI21X1 port map( A => n111, B => n9, C => n71, Y => n174);
   U258 : OAI22X1 port map( A => n112, B => n12, C => n31, D => n114, Y => n175
                           );
   U259 : OAI22X1 port map( A => n114, B => n12, C => n31, D => n211, Y => n176
                           );
   U260 : OAI22X1 port map( A => n211, B => n12, C => n31, D => n212, Y => n177
                           );
   U261 : OAI22X1 port map( A => n212, B => n12, C => n31, D => n213, Y => n178
                           );
   U262 : OAI22X1 port map( A => n213, B => n12, C => n31, D => n214, Y => n179
                           );
   U263 : OAI21X1 port map( A => n214, B => n10, C => n78, Y => n180);
   U264 : OAI22X1 port map( A => n215, B => n11, C => n32, D => n216, Y => n181
                           );
   U265 : OAI22X1 port map( A => n216, B => n11, C => n32, D => n217, Y => n182
                           );
   U266 : OAI22X1 port map( A => n217, B => n11, C => n32, D => n218, Y => n183
                           );
   U267 : OAI22X1 port map( A => n218, B => n12, C => n32, D => n219, Y => n184
                           );
   U268 : OAI22X1 port map( A => n219, B => n11, C => n32, D => n220, Y => n185
                           );
   U269 : OAI21X1 port map( A => n220, B => n10, C => n85, Y => n186);
   U270 : OAI22X1 port map( A => n221, B => n12, C => n32, D => n222, Y => n187
                           );
   U271 : OAI22X1 port map( A => n222, B => n11, C => n32, D => n223, Y => n188
                           );
   U272 : OAI22X1 port map( A => n223, B => n11, C => n33, D => n224, Y => n189
                           );
   U273 : OAI22X1 port map( A => n224, B => n11, C => n33, D => n225, Y => n190
                           );
   U274 : OAI22X1 port map( A => n225, B => n11, C => n33, D => n226, Y => n191
                           );
   U275 : OAI21X1 port map( A => n226, B => n9, C => n92, Y => n192);
   U276 : OAI22X1 port map( A => n227, B => n11, C => n33, D => n228, Y => n193
                           );
   U277 : OAI22X1 port map( A => n228, B => n11, C => n33, D => n229, Y => n194
                           );
   U278 : OAI22X1 port map( A => n229, B => n11, C => n33, D => n230, Y => n195
                           );
   U279 : OAI22X1 port map( A => n230, B => n10, C => n33, D => n231, Y => n196
                           );
   U280 : OAI22X1 port map( A => n231, B => n11, C => n34, D => n232, Y => n197
                           );
   U281 : OAI21X1 port map( A => n232, B => n9, C => n99, Y => n198);
   U282 : OAI22X1 port map( A => n233, B => n10, C => n34, D => n234, Y => n199
                           );
   U283 : OAI22X1 port map( A => n234, B => n10, C => n34, D => n235, Y => n200
                           );
   U284 : OAI22X1 port map( A => n235, B => n10, C => n34, D => n236, Y => n201
                           );
   U285 : OAI22X1 port map( A => n236, B => n10, C => n34, D => n237, Y => n202
                           );
   U286 : OAI22X1 port map( A => n237, B => n10, C => n34, D => n238, Y => n203
                           );
   U287 : OAI21X1 port map( A => n238, B => n9, C => n106, Y => n204);
   U288 : OAI22X1 port map( A => n239, B => n10, C => n34, D => n240, Y => n205
                           );
   U289 : OAI22X1 port map( A => n240, B => n10, C => n35, D => n241, Y => n206
                           );
   U290 : OAI22X1 port map( A => n241, B => n11, C => n35, D => n242, Y => n207
                           );
   U291 : OAI22X1 port map( A => n242, B => n10, C => n35, D => n243, Y => n208
                           );
   U292 : OAI22X1 port map( A => n243, B => n12, C => n35, D => n244, Y => n209
                           );
   U293 : OAI21X1 port map( A => n244, B => n9, C => n113, Y => n210);

end SYN_behavorial;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity world_matrix_buffer is

   port( strb_matrix : in std_logic;  databus_out : in std_logic_vector (15 
         downto 0);  clk : in std_logic;  row_sel : in std_logic_vector (1 
         downto 0);  row : out std_logic_vector (63 downto 0));

end world_matrix_buffer;

architecture SYN_behavorial of world_matrix_buffer is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal regg_255_port, regg_254_port, regg_253_port, regg_252_port, 
      regg_251_port, regg_250_port, regg_249_port, regg_248_port, regg_247_port
      , regg_246_port, regg_245_port, regg_244_port, regg_243_port, 
      regg_242_port, regg_241_port, regg_240_port, regg_239_port, regg_238_port
      , regg_237_port, regg_236_port, regg_235_port, regg_234_port, 
      regg_233_port, regg_232_port, regg_231_port, regg_230_port, regg_229_port
      , regg_228_port, regg_227_port, regg_226_port, regg_225_port, 
      regg_224_port, regg_223_port, regg_222_port, regg_221_port, regg_220_port
      , regg_219_port, regg_218_port, regg_217_port, regg_216_port, 
      regg_215_port, regg_214_port, regg_213_port, regg_212_port, regg_211_port
      , regg_210_port, regg_209_port, regg_208_port, regg_207_port, 
      regg_206_port, regg_205_port, regg_204_port, regg_203_port, regg_202_port
      , regg_201_port, regg_200_port, regg_199_port, regg_198_port, 
      regg_197_port, regg_196_port, regg_195_port, regg_194_port, regg_193_port
      , regg_192_port, regg_191_port, regg_190_port, regg_189_port, 
      regg_188_port, regg_187_port, regg_186_port, regg_185_port, regg_184_port
      , regg_183_port, regg_182_port, regg_181_port, regg_180_port, 
      regg_179_port, regg_178_port, regg_177_port, regg_176_port, regg_175_port
      , regg_174_port, regg_173_port, regg_172_port, regg_171_port, 
      regg_170_port, regg_169_port, regg_168_port, regg_167_port, regg_166_port
      , regg_165_port, regg_164_port, regg_163_port, regg_162_port, 
      regg_161_port, regg_160_port, regg_159_port, regg_158_port, regg_157_port
      , regg_156_port, regg_155_port, regg_154_port, regg_153_port, 
      regg_152_port, regg_151_port, regg_150_port, regg_149_port, regg_148_port
      , regg_147_port, regg_146_port, regg_145_port, regg_144_port, 
      regg_143_port, regg_142_port, regg_141_port, regg_140_port, regg_139_port
      , regg_138_port, regg_137_port, regg_136_port, regg_135_port, 
      regg_134_port, regg_133_port, regg_132_port, regg_131_port, regg_130_port
      , regg_129_port, regg_128_port, regg_127_port, regg_126_port, 
      regg_125_port, regg_124_port, regg_123_port, regg_122_port, regg_121_port
      , regg_120_port, regg_119_port, regg_118_port, regg_117_port, 
      regg_116_port, regg_115_port, regg_114_port, regg_113_port, regg_112_port
      , regg_111_port, regg_110_port, regg_109_port, regg_108_port, 
      regg_107_port, regg_106_port, regg_105_port, regg_104_port, regg_103_port
      , regg_102_port, regg_101_port, regg_100_port, regg_99_port, regg_98_port
      , regg_97_port, regg_96_port, regg_95_port, regg_94_port, regg_93_port, 
      regg_92_port, regg_91_port, regg_90_port, regg_89_port, regg_88_port, 
      regg_87_port, regg_86_port, regg_85_port, regg_84_port, regg_83_port, 
      regg_82_port, regg_81_port, regg_80_port, regg_79_port, regg_78_port, 
      regg_77_port, regg_76_port, regg_75_port, regg_74_port, regg_73_port, 
      regg_72_port, regg_71_port, regg_70_port, regg_69_port, regg_68_port, 
      regg_67_port, regg_66_port, regg_65_port, regg_64_port, regg_63_port, 
      regg_62_port, regg_61_port, regg_60_port, regg_59_port, regg_58_port, 
      regg_57_port, regg_56_port, regg_55_port, regg_54_port, regg_53_port, 
      regg_52_port, regg_51_port, regg_50_port, regg_49_port, regg_48_port, 
      regg_47_port, regg_46_port, regg_45_port, regg_44_port, regg_43_port, 
      regg_42_port, regg_41_port, regg_40_port, regg_39_port, regg_38_port, 
      regg_37_port, regg_36_port, regg_35_port, regg_34_port, regg_33_port, 
      regg_32_port, regg_31_port, regg_30_port, regg_29_port, regg_28_port, 
      regg_27_port, regg_26_port, regg_25_port, regg_24_port, regg_23_port, 
      regg_22_port, regg_21_port, regg_20_port, regg_19_port, regg_18_port, 
      regg_17_port, regg_16_port, regg_15_port, regg_14_port, regg_13_port, 
      regg_12_port, regg_11_port, regg_10_port, regg_9_port, regg_8_port, 
      regg_7_port, regg_6_port, regg_5_port, regg_4_port, regg_3_port, 
      regg_2_port, regg_1_port, regg_0_port, n134, n136, n137, n138, n139, n140
      , n141, n142, n143, n144, n145, n146, n147, n151, n152, n153, n154, n155,
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
      n315, n316, n317, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346, n347, n348, n349, n350, n351, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n372, n373, n374, 
      n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n406, n420, n421, n422, n436, n437, n438, n452, n453, n454, n468, 
      n469, n470, n484, n485, n486, n500, n501, n502, n516, n517, n518, n532, 
      n533, n534, n548, n549, n550, n564, n565, n566, n580, n581, n582, n596, 
      n597, n598, n612, n613, n614, n628, n629, n630, n644, n645, n646, n660, 
      n661, n662, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n135, n148, n149, n150, 
      n165, n166, n167, n182, n183, n184, n199, n200, n201, n216, n217, n218, 
      n233, n234, n235, n250, n251, n252, n267, n268, n269, n284, n285, n286, 
      n301, n302, n303, n318, n319, n320, n335, n336, n337, n352, n353, n354, 
      n369, n370, n371, n386, n387, n388, n403, n404, n405, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, 
      n467, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n583, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
      n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
      n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, 
      n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
      n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, 
      n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, 
      n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, 
      n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, 
      n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804 : 
      std_logic;

begin
   
   regg_reg_15_inst : DFFPOSX1 port map( D => n662, CLK => clk, Q => 
                           regg_15_port);
   regg_reg_31_inst : DFFPOSX1 port map( D => n661, CLK => clk, Q => 
                           regg_31_port);
   regg_reg_47_inst : DFFPOSX1 port map( D => n660, CLK => clk, Q => 
                           regg_47_port);
   regg_reg_63_inst : DFFPOSX1 port map( D => n756, CLK => clk, Q => 
                           regg_63_port);
   regg_reg_79_inst : DFFPOSX1 port map( D => n755, CLK => clk, Q => 
                           regg_79_port);
   regg_reg_95_inst : DFFPOSX1 port map( D => n754, CLK => clk, Q => 
                           regg_95_port);
   regg_reg_111_inst : DFFPOSX1 port map( D => n753, CLK => clk, Q => 
                           regg_111_port);
   regg_reg_127_inst : DFFPOSX1 port map( D => n752, CLK => clk, Q => 
                           regg_127_port);
   regg_reg_143_inst : DFFPOSX1 port map( D => n751, CLK => clk, Q => 
                           regg_143_port);
   regg_reg_159_inst : DFFPOSX1 port map( D => n750, CLK => clk, Q => 
                           regg_159_port);
   regg_reg_175_inst : DFFPOSX1 port map( D => n749, CLK => clk, Q => 
                           regg_175_port);
   regg_reg_191_inst : DFFPOSX1 port map( D => n748, CLK => clk, Q => 
                           regg_191_port);
   regg_reg_207_inst : DFFPOSX1 port map( D => n747, CLK => clk, Q => 
                           regg_207_port);
   regg_reg_223_inst : DFFPOSX1 port map( D => n746, CLK => clk, Q => 
                           regg_223_port);
   regg_reg_239_inst : DFFPOSX1 port map( D => n745, CLK => clk, Q => 
                           regg_239_port);
   regg_reg_255_inst : DFFPOSX1 port map( D => n744, CLK => clk, Q => 
                           regg_255_port);
   regg_reg_14_inst : DFFPOSX1 port map( D => n646, CLK => clk, Q => 
                           regg_14_port);
   regg_reg_30_inst : DFFPOSX1 port map( D => n645, CLK => clk, Q => 
                           regg_30_port);
   regg_reg_46_inst : DFFPOSX1 port map( D => n644, CLK => clk, Q => 
                           regg_46_port);
   regg_reg_62_inst : DFFPOSX1 port map( D => n743, CLK => clk, Q => 
                           regg_62_port);
   regg_reg_78_inst : DFFPOSX1 port map( D => n742, CLK => clk, Q => 
                           regg_78_port);
   regg_reg_94_inst : DFFPOSX1 port map( D => n741, CLK => clk, Q => 
                           regg_94_port);
   regg_reg_110_inst : DFFPOSX1 port map( D => n740, CLK => clk, Q => 
                           regg_110_port);
   regg_reg_126_inst : DFFPOSX1 port map( D => n739, CLK => clk, Q => 
                           regg_126_port);
   regg_reg_142_inst : DFFPOSX1 port map( D => n738, CLK => clk, Q => 
                           regg_142_port);
   regg_reg_158_inst : DFFPOSX1 port map( D => n737, CLK => clk, Q => 
                           regg_158_port);
   regg_reg_174_inst : DFFPOSX1 port map( D => n736, CLK => clk, Q => 
                           regg_174_port);
   regg_reg_190_inst : DFFPOSX1 port map( D => n735, CLK => clk, Q => 
                           regg_190_port);
   regg_reg_206_inst : DFFPOSX1 port map( D => n734, CLK => clk, Q => 
                           regg_206_port);
   regg_reg_222_inst : DFFPOSX1 port map( D => n733, CLK => clk, Q => 
                           regg_222_port);
   regg_reg_238_inst : DFFPOSX1 port map( D => n732, CLK => clk, Q => 
                           regg_238_port);
   regg_reg_254_inst : DFFPOSX1 port map( D => n731, CLK => clk, Q => 
                           regg_254_port);
   regg_reg_13_inst : DFFPOSX1 port map( D => n630, CLK => clk, Q => 
                           regg_13_port);
   regg_reg_29_inst : DFFPOSX1 port map( D => n629, CLK => clk, Q => 
                           regg_29_port);
   regg_reg_45_inst : DFFPOSX1 port map( D => n628, CLK => clk, Q => 
                           regg_45_port);
   regg_reg_61_inst : DFFPOSX1 port map( D => n730, CLK => clk, Q => 
                           regg_61_port);
   regg_reg_77_inst : DFFPOSX1 port map( D => n729, CLK => clk, Q => 
                           regg_77_port);
   regg_reg_93_inst : DFFPOSX1 port map( D => n728, CLK => clk, Q => 
                           regg_93_port);
   regg_reg_109_inst : DFFPOSX1 port map( D => n727, CLK => clk, Q => 
                           regg_109_port);
   regg_reg_125_inst : DFFPOSX1 port map( D => n726, CLK => clk, Q => 
                           regg_125_port);
   regg_reg_141_inst : DFFPOSX1 port map( D => n725, CLK => clk, Q => 
                           regg_141_port);
   regg_reg_157_inst : DFFPOSX1 port map( D => n724, CLK => clk, Q => 
                           regg_157_port);
   regg_reg_173_inst : DFFPOSX1 port map( D => n723, CLK => clk, Q => 
                           regg_173_port);
   regg_reg_189_inst : DFFPOSX1 port map( D => n722, CLK => clk, Q => 
                           regg_189_port);
   regg_reg_205_inst : DFFPOSX1 port map( D => n721, CLK => clk, Q => 
                           regg_205_port);
   regg_reg_221_inst : DFFPOSX1 port map( D => n720, CLK => clk, Q => 
                           regg_221_port);
   regg_reg_237_inst : DFFPOSX1 port map( D => n719, CLK => clk, Q => 
                           regg_237_port);
   regg_reg_253_inst : DFFPOSX1 port map( D => n718, CLK => clk, Q => 
                           regg_253_port);
   regg_reg_12_inst : DFFPOSX1 port map( D => n614, CLK => clk, Q => 
                           regg_12_port);
   regg_reg_28_inst : DFFPOSX1 port map( D => n613, CLK => clk, Q => 
                           regg_28_port);
   regg_reg_44_inst : DFFPOSX1 port map( D => n612, CLK => clk, Q => 
                           regg_44_port);
   regg_reg_60_inst : DFFPOSX1 port map( D => n717, CLK => clk, Q => 
                           regg_60_port);
   regg_reg_76_inst : DFFPOSX1 port map( D => n716, CLK => clk, Q => 
                           regg_76_port);
   regg_reg_92_inst : DFFPOSX1 port map( D => n715, CLK => clk, Q => 
                           regg_92_port);
   regg_reg_108_inst : DFFPOSX1 port map( D => n714, CLK => clk, Q => 
                           regg_108_port);
   regg_reg_124_inst : DFFPOSX1 port map( D => n713, CLK => clk, Q => 
                           regg_124_port);
   regg_reg_140_inst : DFFPOSX1 port map( D => n712, CLK => clk, Q => 
                           regg_140_port);
   regg_reg_156_inst : DFFPOSX1 port map( D => n711, CLK => clk, Q => 
                           regg_156_port);
   regg_reg_172_inst : DFFPOSX1 port map( D => n710, CLK => clk, Q => 
                           regg_172_port);
   regg_reg_188_inst : DFFPOSX1 port map( D => n709, CLK => clk, Q => 
                           regg_188_port);
   regg_reg_204_inst : DFFPOSX1 port map( D => n708, CLK => clk, Q => 
                           regg_204_port);
   regg_reg_220_inst : DFFPOSX1 port map( D => n707, CLK => clk, Q => 
                           regg_220_port);
   regg_reg_236_inst : DFFPOSX1 port map( D => n706, CLK => clk, Q => 
                           regg_236_port);
   regg_reg_252_inst : DFFPOSX1 port map( D => n705, CLK => clk, Q => 
                           regg_252_port);
   regg_reg_11_inst : DFFPOSX1 port map( D => n598, CLK => clk, Q => 
                           regg_11_port);
   regg_reg_27_inst : DFFPOSX1 port map( D => n597, CLK => clk, Q => 
                           regg_27_port);
   regg_reg_43_inst : DFFPOSX1 port map( D => n596, CLK => clk, Q => 
                           regg_43_port);
   regg_reg_59_inst : DFFPOSX1 port map( D => n704, CLK => clk, Q => 
                           regg_59_port);
   regg_reg_75_inst : DFFPOSX1 port map( D => n703, CLK => clk, Q => 
                           regg_75_port);
   regg_reg_91_inst : DFFPOSX1 port map( D => n702, CLK => clk, Q => 
                           regg_91_port);
   regg_reg_107_inst : DFFPOSX1 port map( D => n701, CLK => clk, Q => 
                           regg_107_port);
   regg_reg_123_inst : DFFPOSX1 port map( D => n700, CLK => clk, Q => 
                           regg_123_port);
   regg_reg_139_inst : DFFPOSX1 port map( D => n699, CLK => clk, Q => 
                           regg_139_port);
   regg_reg_155_inst : DFFPOSX1 port map( D => n698, CLK => clk, Q => 
                           regg_155_port);
   regg_reg_171_inst : DFFPOSX1 port map( D => n697, CLK => clk, Q => 
                           regg_171_port);
   regg_reg_187_inst : DFFPOSX1 port map( D => n696, CLK => clk, Q => 
                           regg_187_port);
   regg_reg_203_inst : DFFPOSX1 port map( D => n695, CLK => clk, Q => 
                           regg_203_port);
   regg_reg_219_inst : DFFPOSX1 port map( D => n694, CLK => clk, Q => 
                           regg_219_port);
   regg_reg_235_inst : DFFPOSX1 port map( D => n693, CLK => clk, Q => 
                           regg_235_port);
   regg_reg_251_inst : DFFPOSX1 port map( D => n692, CLK => clk, Q => 
                           regg_251_port);
   regg_reg_10_inst : DFFPOSX1 port map( D => n582, CLK => clk, Q => 
                           regg_10_port);
   regg_reg_26_inst : DFFPOSX1 port map( D => n581, CLK => clk, Q => 
                           regg_26_port);
   regg_reg_42_inst : DFFPOSX1 port map( D => n580, CLK => clk, Q => 
                           regg_42_port);
   regg_reg_58_inst : DFFPOSX1 port map( D => n691, CLK => clk, Q => 
                           regg_58_port);
   regg_reg_74_inst : DFFPOSX1 port map( D => n690, CLK => clk, Q => 
                           regg_74_port);
   regg_reg_90_inst : DFFPOSX1 port map( D => n689, CLK => clk, Q => 
                           regg_90_port);
   regg_reg_106_inst : DFFPOSX1 port map( D => n688, CLK => clk, Q => 
                           regg_106_port);
   regg_reg_122_inst : DFFPOSX1 port map( D => n687, CLK => clk, Q => 
                           regg_122_port);
   regg_reg_138_inst : DFFPOSX1 port map( D => n686, CLK => clk, Q => 
                           regg_138_port);
   regg_reg_154_inst : DFFPOSX1 port map( D => n685, CLK => clk, Q => 
                           regg_154_port);
   regg_reg_170_inst : DFFPOSX1 port map( D => n684, CLK => clk, Q => 
                           regg_170_port);
   regg_reg_186_inst : DFFPOSX1 port map( D => n683, CLK => clk, Q => 
                           regg_186_port);
   regg_reg_202_inst : DFFPOSX1 port map( D => n682, CLK => clk, Q => 
                           regg_202_port);
   regg_reg_218_inst : DFFPOSX1 port map( D => n681, CLK => clk, Q => 
                           regg_218_port);
   regg_reg_234_inst : DFFPOSX1 port map( D => n680, CLK => clk, Q => 
                           regg_234_port);
   regg_reg_250_inst : DFFPOSX1 port map( D => n679, CLK => clk, Q => 
                           regg_250_port);
   regg_reg_9_inst : DFFPOSX1 port map( D => n566, CLK => clk, Q => regg_9_port
                           );
   regg_reg_25_inst : DFFPOSX1 port map( D => n565, CLK => clk, Q => 
                           regg_25_port);
   regg_reg_41_inst : DFFPOSX1 port map( D => n564, CLK => clk, Q => 
                           regg_41_port);
   regg_reg_57_inst : DFFPOSX1 port map( D => n678, CLK => clk, Q => 
                           regg_57_port);
   regg_reg_73_inst : DFFPOSX1 port map( D => n677, CLK => clk, Q => 
                           regg_73_port);
   regg_reg_89_inst : DFFPOSX1 port map( D => n676, CLK => clk, Q => 
                           regg_89_port);
   regg_reg_105_inst : DFFPOSX1 port map( D => n675, CLK => clk, Q => 
                           regg_105_port);
   regg_reg_121_inst : DFFPOSX1 port map( D => n674, CLK => clk, Q => 
                           regg_121_port);
   regg_reg_137_inst : DFFPOSX1 port map( D => n673, CLK => clk, Q => 
                           regg_137_port);
   regg_reg_153_inst : DFFPOSX1 port map( D => n672, CLK => clk, Q => 
                           regg_153_port);
   regg_reg_169_inst : DFFPOSX1 port map( D => n671, CLK => clk, Q => 
                           regg_169_port);
   regg_reg_185_inst : DFFPOSX1 port map( D => n670, CLK => clk, Q => 
                           regg_185_port);
   regg_reg_201_inst : DFFPOSX1 port map( D => n669, CLK => clk, Q => 
                           regg_201_port);
   regg_reg_217_inst : DFFPOSX1 port map( D => n668, CLK => clk, Q => 
                           regg_217_port);
   regg_reg_233_inst : DFFPOSX1 port map( D => n667, CLK => clk, Q => 
                           regg_233_port);
   regg_reg_249_inst : DFFPOSX1 port map( D => n666, CLK => clk, Q => 
                           regg_249_port);
   regg_reg_8_inst : DFFPOSX1 port map( D => n550, CLK => clk, Q => regg_8_port
                           );
   regg_reg_24_inst : DFFPOSX1 port map( D => n549, CLK => clk, Q => 
                           regg_24_port);
   regg_reg_40_inst : DFFPOSX1 port map( D => n548, CLK => clk, Q => 
                           regg_40_port);
   regg_reg_56_inst : DFFPOSX1 port map( D => n665, CLK => clk, Q => 
                           regg_56_port);
   regg_reg_72_inst : DFFPOSX1 port map( D => n664, CLK => clk, Q => 
                           regg_72_port);
   regg_reg_88_inst : DFFPOSX1 port map( D => n663, CLK => clk, Q => 
                           regg_88_port);
   regg_reg_104_inst : DFFPOSX1 port map( D => n659, CLK => clk, Q => 
                           regg_104_port);
   regg_reg_120_inst : DFFPOSX1 port map( D => n658, CLK => clk, Q => 
                           regg_120_port);
   regg_reg_136_inst : DFFPOSX1 port map( D => n657, CLK => clk, Q => 
                           regg_136_port);
   regg_reg_152_inst : DFFPOSX1 port map( D => n656, CLK => clk, Q => 
                           regg_152_port);
   regg_reg_168_inst : DFFPOSX1 port map( D => n655, CLK => clk, Q => 
                           regg_168_port);
   regg_reg_184_inst : DFFPOSX1 port map( D => n654, CLK => clk, Q => 
                           regg_184_port);
   regg_reg_200_inst : DFFPOSX1 port map( D => n653, CLK => clk, Q => 
                           regg_200_port);
   regg_reg_216_inst : DFFPOSX1 port map( D => n652, CLK => clk, Q => 
                           regg_216_port);
   regg_reg_232_inst : DFFPOSX1 port map( D => n651, CLK => clk, Q => 
                           regg_232_port);
   regg_reg_248_inst : DFFPOSX1 port map( D => n650, CLK => clk, Q => 
                           regg_248_port);
   regg_reg_7_inst : DFFPOSX1 port map( D => n534, CLK => clk, Q => regg_7_port
                           );
   regg_reg_23_inst : DFFPOSX1 port map( D => n533, CLK => clk, Q => 
                           regg_23_port);
   regg_reg_39_inst : DFFPOSX1 port map( D => n532, CLK => clk, Q => 
                           regg_39_port);
   regg_reg_55_inst : DFFPOSX1 port map( D => n649, CLK => clk, Q => 
                           regg_55_port);
   regg_reg_71_inst : DFFPOSX1 port map( D => n648, CLK => clk, Q => 
                           regg_71_port);
   regg_reg_87_inst : DFFPOSX1 port map( D => n647, CLK => clk, Q => 
                           regg_87_port);
   regg_reg_103_inst : DFFPOSX1 port map( D => n643, CLK => clk, Q => 
                           regg_103_port);
   regg_reg_119_inst : DFFPOSX1 port map( D => n642, CLK => clk, Q => 
                           regg_119_port);
   regg_reg_135_inst : DFFPOSX1 port map( D => n641, CLK => clk, Q => 
                           regg_135_port);
   regg_reg_151_inst : DFFPOSX1 port map( D => n640, CLK => clk, Q => 
                           regg_151_port);
   regg_reg_167_inst : DFFPOSX1 port map( D => n639, CLK => clk, Q => 
                           regg_167_port);
   regg_reg_183_inst : DFFPOSX1 port map( D => n638, CLK => clk, Q => 
                           regg_183_port);
   regg_reg_199_inst : DFFPOSX1 port map( D => n637, CLK => clk, Q => 
                           regg_199_port);
   regg_reg_215_inst : DFFPOSX1 port map( D => n636, CLK => clk, Q => 
                           regg_215_port);
   regg_reg_231_inst : DFFPOSX1 port map( D => n635, CLK => clk, Q => 
                           regg_231_port);
   regg_reg_247_inst : DFFPOSX1 port map( D => n634, CLK => clk, Q => 
                           regg_247_port);
   regg_reg_6_inst : DFFPOSX1 port map( D => n518, CLK => clk, Q => regg_6_port
                           );
   regg_reg_22_inst : DFFPOSX1 port map( D => n517, CLK => clk, Q => 
                           regg_22_port);
   regg_reg_38_inst : DFFPOSX1 port map( D => n516, CLK => clk, Q => 
                           regg_38_port);
   regg_reg_54_inst : DFFPOSX1 port map( D => n633, CLK => clk, Q => 
                           regg_54_port);
   regg_reg_70_inst : DFFPOSX1 port map( D => n632, CLK => clk, Q => 
                           regg_70_port);
   regg_reg_86_inst : DFFPOSX1 port map( D => n631, CLK => clk, Q => 
                           regg_86_port);
   regg_reg_102_inst : DFFPOSX1 port map( D => n627, CLK => clk, Q => 
                           regg_102_port);
   regg_reg_118_inst : DFFPOSX1 port map( D => n626, CLK => clk, Q => 
                           regg_118_port);
   regg_reg_134_inst : DFFPOSX1 port map( D => n625, CLK => clk, Q => 
                           regg_134_port);
   regg_reg_150_inst : DFFPOSX1 port map( D => n624, CLK => clk, Q => 
                           regg_150_port);
   regg_reg_166_inst : DFFPOSX1 port map( D => n623, CLK => clk, Q => 
                           regg_166_port);
   regg_reg_182_inst : DFFPOSX1 port map( D => n622, CLK => clk, Q => 
                           regg_182_port);
   regg_reg_198_inst : DFFPOSX1 port map( D => n621, CLK => clk, Q => 
                           regg_198_port);
   regg_reg_214_inst : DFFPOSX1 port map( D => n620, CLK => clk, Q => 
                           regg_214_port);
   regg_reg_230_inst : DFFPOSX1 port map( D => n619, CLK => clk, Q => 
                           regg_230_port);
   regg_reg_246_inst : DFFPOSX1 port map( D => n618, CLK => clk, Q => 
                           regg_246_port);
   regg_reg_5_inst : DFFPOSX1 port map( D => n502, CLK => clk, Q => regg_5_port
                           );
   regg_reg_21_inst : DFFPOSX1 port map( D => n501, CLK => clk, Q => 
                           regg_21_port);
   regg_reg_37_inst : DFFPOSX1 port map( D => n500, CLK => clk, Q => 
                           regg_37_port);
   regg_reg_53_inst : DFFPOSX1 port map( D => n617, CLK => clk, Q => 
                           regg_53_port);
   regg_reg_69_inst : DFFPOSX1 port map( D => n616, CLK => clk, Q => 
                           regg_69_port);
   regg_reg_85_inst : DFFPOSX1 port map( D => n615, CLK => clk, Q => 
                           regg_85_port);
   regg_reg_101_inst : DFFPOSX1 port map( D => n611, CLK => clk, Q => 
                           regg_101_port);
   regg_reg_117_inst : DFFPOSX1 port map( D => n610, CLK => clk, Q => 
                           regg_117_port);
   regg_reg_133_inst : DFFPOSX1 port map( D => n609, CLK => clk, Q => 
                           regg_133_port);
   regg_reg_149_inst : DFFPOSX1 port map( D => n608, CLK => clk, Q => 
                           regg_149_port);
   regg_reg_165_inst : DFFPOSX1 port map( D => n607, CLK => clk, Q => 
                           regg_165_port);
   regg_reg_181_inst : DFFPOSX1 port map( D => n606, CLK => clk, Q => 
                           regg_181_port);
   regg_reg_197_inst : DFFPOSX1 port map( D => n605, CLK => clk, Q => 
                           regg_197_port);
   regg_reg_213_inst : DFFPOSX1 port map( D => n604, CLK => clk, Q => 
                           regg_213_port);
   regg_reg_229_inst : DFFPOSX1 port map( D => n603, CLK => clk, Q => 
                           regg_229_port);
   regg_reg_245_inst : DFFPOSX1 port map( D => n602, CLK => clk, Q => 
                           regg_245_port);
   regg_reg_4_inst : DFFPOSX1 port map( D => n486, CLK => clk, Q => regg_4_port
                           );
   regg_reg_20_inst : DFFPOSX1 port map( D => n485, CLK => clk, Q => 
                           regg_20_port);
   regg_reg_36_inst : DFFPOSX1 port map( D => n484, CLK => clk, Q => 
                           regg_36_port);
   regg_reg_52_inst : DFFPOSX1 port map( D => n601, CLK => clk, Q => 
                           regg_52_port);
   regg_reg_68_inst : DFFPOSX1 port map( D => n600, CLK => clk, Q => 
                           regg_68_port);
   regg_reg_84_inst : DFFPOSX1 port map( D => n599, CLK => clk, Q => 
                           regg_84_port);
   regg_reg_100_inst : DFFPOSX1 port map( D => n595, CLK => clk, Q => 
                           regg_100_port);
   regg_reg_116_inst : DFFPOSX1 port map( D => n594, CLK => clk, Q => 
                           regg_116_port);
   regg_reg_132_inst : DFFPOSX1 port map( D => n593, CLK => clk, Q => 
                           regg_132_port);
   regg_reg_148_inst : DFFPOSX1 port map( D => n592, CLK => clk, Q => 
                           regg_148_port);
   regg_reg_164_inst : DFFPOSX1 port map( D => n591, CLK => clk, Q => 
                           regg_164_port);
   regg_reg_180_inst : DFFPOSX1 port map( D => n590, CLK => clk, Q => 
                           regg_180_port);
   regg_reg_196_inst : DFFPOSX1 port map( D => n589, CLK => clk, Q => 
                           regg_196_port);
   regg_reg_212_inst : DFFPOSX1 port map( D => n588, CLK => clk, Q => 
                           regg_212_port);
   regg_reg_228_inst : DFFPOSX1 port map( D => n587, CLK => clk, Q => 
                           regg_228_port);
   regg_reg_244_inst : DFFPOSX1 port map( D => n586, CLK => clk, Q => 
                           regg_244_port);
   regg_reg_3_inst : DFFPOSX1 port map( D => n470, CLK => clk, Q => regg_3_port
                           );
   regg_reg_19_inst : DFFPOSX1 port map( D => n469, CLK => clk, Q => 
                           regg_19_port);
   regg_reg_35_inst : DFFPOSX1 port map( D => n468, CLK => clk, Q => 
                           regg_35_port);
   regg_reg_51_inst : DFFPOSX1 port map( D => n585, CLK => clk, Q => 
                           regg_51_port);
   regg_reg_67_inst : DFFPOSX1 port map( D => n584, CLK => clk, Q => 
                           regg_67_port);
   regg_reg_83_inst : DFFPOSX1 port map( D => n583, CLK => clk, Q => 
                           regg_83_port);
   regg_reg_99_inst : DFFPOSX1 port map( D => n579, CLK => clk, Q => 
                           regg_99_port);
   regg_reg_115_inst : DFFPOSX1 port map( D => n578, CLK => clk, Q => 
                           regg_115_port);
   regg_reg_131_inst : DFFPOSX1 port map( D => n577, CLK => clk, Q => 
                           regg_131_port);
   regg_reg_147_inst : DFFPOSX1 port map( D => n576, CLK => clk, Q => 
                           regg_147_port);
   regg_reg_163_inst : DFFPOSX1 port map( D => n575, CLK => clk, Q => 
                           regg_163_port);
   regg_reg_179_inst : DFFPOSX1 port map( D => n574, CLK => clk, Q => 
                           regg_179_port);
   regg_reg_195_inst : DFFPOSX1 port map( D => n573, CLK => clk, Q => 
                           regg_195_port);
   regg_reg_211_inst : DFFPOSX1 port map( D => n572, CLK => clk, Q => 
                           regg_211_port);
   regg_reg_227_inst : DFFPOSX1 port map( D => n571, CLK => clk, Q => 
                           regg_227_port);
   regg_reg_243_inst : DFFPOSX1 port map( D => n570, CLK => clk, Q => 
                           regg_243_port);
   regg_reg_2_inst : DFFPOSX1 port map( D => n454, CLK => clk, Q => regg_2_port
                           );
   regg_reg_18_inst : DFFPOSX1 port map( D => n453, CLK => clk, Q => 
                           regg_18_port);
   regg_reg_34_inst : DFFPOSX1 port map( D => n452, CLK => clk, Q => 
                           regg_34_port);
   regg_reg_50_inst : DFFPOSX1 port map( D => n569, CLK => clk, Q => 
                           regg_50_port);
   regg_reg_66_inst : DFFPOSX1 port map( D => n568, CLK => clk, Q => 
                           regg_66_port);
   regg_reg_82_inst : DFFPOSX1 port map( D => n567, CLK => clk, Q => 
                           regg_82_port);
   regg_reg_98_inst : DFFPOSX1 port map( D => n563, CLK => clk, Q => 
                           regg_98_port);
   regg_reg_114_inst : DFFPOSX1 port map( D => n562, CLK => clk, Q => 
                           regg_114_port);
   regg_reg_130_inst : DFFPOSX1 port map( D => n561, CLK => clk, Q => 
                           regg_130_port);
   regg_reg_146_inst : DFFPOSX1 port map( D => n560, CLK => clk, Q => 
                           regg_146_port);
   regg_reg_162_inst : DFFPOSX1 port map( D => n559, CLK => clk, Q => 
                           regg_162_port);
   regg_reg_178_inst : DFFPOSX1 port map( D => n558, CLK => clk, Q => 
                           regg_178_port);
   regg_reg_194_inst : DFFPOSX1 port map( D => n557, CLK => clk, Q => 
                           regg_194_port);
   regg_reg_210_inst : DFFPOSX1 port map( D => n556, CLK => clk, Q => 
                           regg_210_port);
   regg_reg_226_inst : DFFPOSX1 port map( D => n555, CLK => clk, Q => 
                           regg_226_port);
   regg_reg_242_inst : DFFPOSX1 port map( D => n554, CLK => clk, Q => 
                           regg_242_port);
   regg_reg_1_inst : DFFPOSX1 port map( D => n438, CLK => clk, Q => regg_1_port
                           );
   regg_reg_17_inst : DFFPOSX1 port map( D => n437, CLK => clk, Q => 
                           regg_17_port);
   regg_reg_33_inst : DFFPOSX1 port map( D => n436, CLK => clk, Q => 
                           regg_33_port);
   regg_reg_49_inst : DFFPOSX1 port map( D => n553, CLK => clk, Q => 
                           regg_49_port);
   regg_reg_65_inst : DFFPOSX1 port map( D => n552, CLK => clk, Q => 
                           regg_65_port);
   regg_reg_81_inst : DFFPOSX1 port map( D => n551, CLK => clk, Q => 
                           regg_81_port);
   regg_reg_97_inst : DFFPOSX1 port map( D => n547, CLK => clk, Q => 
                           regg_97_port);
   regg_reg_113_inst : DFFPOSX1 port map( D => n546, CLK => clk, Q => 
                           regg_113_port);
   regg_reg_129_inst : DFFPOSX1 port map( D => n545, CLK => clk, Q => 
                           regg_129_port);
   regg_reg_145_inst : DFFPOSX1 port map( D => n544, CLK => clk, Q => 
                           regg_145_port);
   regg_reg_161_inst : DFFPOSX1 port map( D => n543, CLK => clk, Q => 
                           regg_161_port);
   regg_reg_177_inst : DFFPOSX1 port map( D => n542, CLK => clk, Q => 
                           regg_177_port);
   regg_reg_193_inst : DFFPOSX1 port map( D => n541, CLK => clk, Q => 
                           regg_193_port);
   regg_reg_209_inst : DFFPOSX1 port map( D => n540, CLK => clk, Q => 
                           regg_209_port);
   regg_reg_225_inst : DFFPOSX1 port map( D => n539, CLK => clk, Q => 
                           regg_225_port);
   regg_reg_241_inst : DFFPOSX1 port map( D => n538, CLK => clk, Q => 
                           regg_241_port);
   regg_reg_0_inst : DFFPOSX1 port map( D => n422, CLK => clk, Q => regg_0_port
                           );
   regg_reg_16_inst : DFFPOSX1 port map( D => n421, CLK => clk, Q => 
                           regg_16_port);
   regg_reg_32_inst : DFFPOSX1 port map( D => n420, CLK => clk, Q => 
                           regg_32_port);
   regg_reg_48_inst : DFFPOSX1 port map( D => n537, CLK => clk, Q => 
                           regg_48_port);
   regg_reg_64_inst : DFFPOSX1 port map( D => n536, CLK => clk, Q => 
                           regg_64_port);
   regg_reg_80_inst : DFFPOSX1 port map( D => n535, CLK => clk, Q => 
                           regg_80_port);
   regg_reg_96_inst : DFFPOSX1 port map( D => n531, CLK => clk, Q => 
                           regg_96_port);
   regg_reg_112_inst : DFFPOSX1 port map( D => n530, CLK => clk, Q => 
                           regg_112_port);
   regg_reg_128_inst : DFFPOSX1 port map( D => n529, CLK => clk, Q => 
                           regg_128_port);
   regg_reg_144_inst : DFFPOSX1 port map( D => n528, CLK => clk, Q => 
                           regg_144_port);
   regg_reg_160_inst : DFFPOSX1 port map( D => n527, CLK => clk, Q => 
                           regg_160_port);
   regg_reg_176_inst : DFFPOSX1 port map( D => n526, CLK => clk, Q => 
                           regg_176_port);
   regg_reg_192_inst : DFFPOSX1 port map( D => n525, CLK => clk, Q => 
                           regg_192_port);
   regg_reg_208_inst : DFFPOSX1 port map( D => n524, CLK => clk, Q => 
                           regg_208_port);
   regg_reg_224_inst : DFFPOSX1 port map( D => n523, CLK => clk, Q => 
                           regg_224_port);
   regg_reg_240_inst : DFFPOSX1 port map( D => n522, CLK => clk, Q => 
                           regg_240_port);
   U200 : AOI22X1 port map( A => n96, B => regg_240_port, C => regg_224_port, D
                           => n46, Y => n134);
   U202 : AOI22X1 port map( A => n96, B => regg_224_port, C => regg_208_port, D
                           => n46, Y => n136);
   U204 : AOI22X1 port map( A => n96, B => regg_208_port, C => regg_192_port, D
                           => n46, Y => n137);
   U206 : AOI22X1 port map( A => n95, B => regg_192_port, C => regg_176_port, D
                           => n46, Y => n138);
   U208 : AOI22X1 port map( A => n95, B => regg_176_port, C => regg_160_port, D
                           => n47, Y => n139);
   U210 : AOI22X1 port map( A => n94, B => regg_160_port, C => regg_144_port, D
                           => n47, Y => n140);
   U212 : AOI22X1 port map( A => n94, B => regg_144_port, C => regg_128_port, D
                           => n47, Y => n141);
   U214 : AOI22X1 port map( A => n92, B => regg_128_port, C => regg_112_port, D
                           => n47, Y => n142);
   U216 : AOI22X1 port map( A => regg_96_port, B => n60, C => n75, D => 
                           regg_112_port, Y => n143);
   U218 : AOI22X1 port map( A => n92, B => regg_96_port, C => regg_80_port, D 
                           => n47, Y => n144);
   U220 : AOI22X1 port map( A => n92, B => regg_80_port, C => regg_64_port, D 
                           => n47, Y => n145);
   U222 : AOI22X1 port map( A => n91, B => regg_64_port, C => regg_48_port, D 
                           => n46, Y => n146);
   U224 : AOI22X1 port map( A => n91, B => regg_48_port, C => regg_32_port, D 
                           => n46, Y => n147);
   U225 : OAI22X1 port map( A => n62, B => n804, C => n803, D => n73, Y => n420
                           );
   U227 : OAI22X1 port map( A => n62, B => n803, C => n802, D => n71, Y => n421
                           );
   U229 : OAI21X1 port map( A => n65, B => n802, C => n151, Y => n422);
   U230 : NAND2X1 port map( A => databus_out(0), B => n64, Y => n151);
   U233 : AOI22X1 port map( A => n91, B => regg_241_port, C => regg_225_port, D
                           => n47, Y => n152);
   U235 : AOI22X1 port map( A => n89, B => regg_225_port, C => regg_209_port, D
                           => n57, Y => n153);
   U237 : AOI22X1 port map( A => n88, B => regg_209_port, C => regg_193_port, D
                           => n48, Y => n154);
   U239 : AOI22X1 port map( A => n88, B => regg_193_port, C => regg_177_port, D
                           => n48, Y => n155);
   U241 : AOI22X1 port map( A => n88, B => regg_177_port, C => regg_161_port, D
                           => n48, Y => n156);
   U243 : AOI22X1 port map( A => n87, B => regg_161_port, C => regg_145_port, D
                           => n48, Y => n157);
   U245 : AOI22X1 port map( A => n86, B => regg_145_port, C => regg_129_port, D
                           => n48, Y => n158);
   U247 : AOI22X1 port map( A => n85, B => regg_129_port, C => regg_113_port, D
                           => n48, Y => n159);
   U249 : AOI22X1 port map( A => regg_97_port, B => n60, C => n77, D => 
                           regg_113_port, Y => n160);
   U251 : AOI22X1 port map( A => n85, B => regg_97_port, C => regg_81_port, D 
                           => n57, Y => n161);
   U253 : AOI22X1 port map( A => n85, B => regg_81_port, C => regg_65_port, D 
                           => n48, Y => n162);
   U255 : AOI22X1 port map( A => n84, B => regg_65_port, C => regg_49_port, D 
                           => n57, Y => n163);
   U257 : AOI22X1 port map( A => n83, B => regg_49_port, C => regg_33_port, D 
                           => n58, Y => n164);
   U258 : OAI22X1 port map( A => n64, B => n801, C => n800, D => n73, Y => n436
                           );
   U260 : OAI22X1 port map( A => n799, B => n79, C => n62, D => n800, Y => n437
                           );
   U262 : OAI21X1 port map( A => n64, B => n799, C => n168, Y => n438);
   U263 : NAND2X1 port map( A => databus_out(1), B => n65, Y => n168);
   U266 : AOI22X1 port map( A => n82, B => regg_242_port, C => regg_226_port, D
                           => n49, Y => n169);
   U268 : AOI22X1 port map( A => n82, B => regg_226_port, C => regg_210_port, D
                           => n49, Y => n170);
   U270 : AOI22X1 port map( A => n81, B => regg_210_port, C => regg_194_port, D
                           => n58, Y => n171);
   U272 : AOI22X1 port map( A => n81, B => regg_194_port, C => regg_178_port, D
                           => n49, Y => n172);
   U274 : AOI22X1 port map( A => n80, B => regg_178_port, C => regg_162_port, D
                           => n49, Y => n173);
   U276 : AOI22X1 port map( A => n80, B => regg_162_port, C => regg_146_port, D
                           => n49, Y => n174);
   U278 : AOI22X1 port map( A => n79, B => regg_146_port, C => regg_130_port, D
                           => n49, Y => n175);
   U280 : AOI22X1 port map( A => n80, B => regg_130_port, C => regg_114_port, D
                           => n49, Y => n176);
   U282 : AOI22X1 port map( A => regg_98_port, B => n61, C => n77, D => 
                           regg_114_port, Y => n177);
   U284 : AOI22X1 port map( A => n80, B => regg_98_port, C => regg_82_port, D 
                           => n49, Y => n178);
   U286 : AOI22X1 port map( A => n80, B => regg_82_port, C => regg_66_port, D 
                           => n50, Y => n179);
   U288 : AOI22X1 port map( A => n81, B => regg_66_port, C => regg_50_port, D 
                           => n50, Y => n180);
   U290 : AOI22X1 port map( A => n81, B => regg_50_port, C => regg_34_port, D 
                           => n58, Y => n181);
   U291 : OAI22X1 port map( A => n63, B => n798, C => n797, D => n74, Y => n452
                           );
   U293 : OAI22X1 port map( A => n796, B => n78, C => n62, D => n797, Y => n453
                           );
   U295 : OAI21X1 port map( A => n64, B => n796, C => n185, Y => n454);
   U296 : NAND2X1 port map( A => databus_out(2), B => n65, Y => n185);
   U299 : AOI22X1 port map( A => n81, B => regg_243_port, C => regg_227_port, D
                           => n59, Y => n186);
   U301 : AOI22X1 port map( A => n82, B => regg_227_port, C => regg_211_port, D
                           => n59, Y => n187);
   U303 : AOI22X1 port map( A => n82, B => regg_211_port, C => regg_195_port, D
                           => n50, Y => n188);
   U305 : AOI22X1 port map( A => n82, B => regg_195_port, C => regg_179_port, D
                           => n50, Y => n189);
   U307 : AOI22X1 port map( A => n83, B => regg_179_port, C => regg_163_port, D
                           => n50, Y => n190);
   U309 : AOI22X1 port map( A => n83, B => regg_163_port, C => regg_147_port, D
                           => n59, Y => n191);
   U311 : AOI22X1 port map( A => n83, B => regg_147_port, C => regg_131_port, D
                           => n51, Y => n192);
   U313 : AOI22X1 port map( A => n83, B => regg_131_port, C => regg_115_port, D
                           => n51, Y => n193);
   U315 : AOI22X1 port map( A => regg_99_port, B => n61, C => n76, D => 
                           regg_115_port, Y => n194);
   U317 : AOI22X1 port map( A => n84, B => regg_99_port, C => regg_83_port, D 
                           => n59, Y => n195);
   U319 : AOI22X1 port map( A => n84, B => regg_83_port, C => regg_67_port, D 
                           => n51, Y => n196);
   U321 : AOI22X1 port map( A => n84, B => regg_67_port, C => regg_51_port, D 
                           => n58, Y => n197);
   U323 : AOI22X1 port map( A => n84, B => regg_51_port, C => regg_35_port, D 
                           => n58, Y => n198);
   U324 : OAI22X1 port map( A => n64, B => n795, C => n794, D => n73, Y => n468
                           );
   U326 : OAI22X1 port map( A => n793, B => n79, C => n62, D => n794, Y => n469
                           );
   U328 : OAI21X1 port map( A => n65, B => n793, C => n202, Y => n470);
   U329 : NAND2X1 port map( A => databus_out(3), B => n65, Y => n202);
   U332 : AOI22X1 port map( A => n85, B => regg_244_port, C => regg_228_port, D
                           => n51, Y => n203);
   U334 : AOI22X1 port map( A => n85, B => regg_228_port, C => regg_212_port, D
                           => n51, Y => n204);
   U336 : AOI22X1 port map( A => n86, B => regg_212_port, C => regg_196_port, D
                           => n51, Y => n205);
   U338 : AOI22X1 port map( A => n86, B => regg_196_port, C => regg_180_port, D
                           => n52, Y => n206);
   U340 : AOI22X1 port map( A => n86, B => regg_180_port, C => regg_164_port, D
                           => n57, Y => n207);
   U342 : AOI22X1 port map( A => n86, B => regg_164_port, C => regg_148_port, D
                           => n52, Y => n208);
   U344 : AOI22X1 port map( A => n87, B => regg_148_port, C => regg_132_port, D
                           => n52, Y => n209);
   U346 : AOI22X1 port map( A => n87, B => regg_132_port, C => regg_116_port, D
                           => n52, Y => n210);
   U348 : AOI22X1 port map( A => n87, B => regg_116_port, C => regg_100_port, D
                           => n52, Y => n211);
   U350 : AOI22X1 port map( A => regg_84_port, B => n61, C => n76, D => 
                           regg_100_port, Y => n212);
   U352 : AOI22X1 port map( A => n87, B => regg_84_port, C => regg_68_port, D 
                           => n52, Y => n213);
   U354 : AOI22X1 port map( A => n88, B => regg_68_port, C => regg_52_port, D 
                           => n56, Y => n214);
   U356 : AOI22X1 port map( A => n88, B => regg_52_port, C => regg_36_port, D 
                           => n56, Y => n215);
   U357 : OAI22X1 port map( A => n63, B => n792, C => n791, D => n73, Y => n484
                           );
   U359 : OAI22X1 port map( A => n790, B => n79, C => n62, D => n791, Y => n485
                           );
   U361 : OAI21X1 port map( A => n65, B => n790, C => n219, Y => n486);
   U362 : NAND2X1 port map( A => databus_out(4), B => n63, Y => n219);
   U365 : AOI22X1 port map( A => n89, B => regg_245_port, C => regg_229_port, D
                           => n52, Y => n220);
   U367 : AOI22X1 port map( A => n89, B => regg_229_port, C => regg_213_port, D
                           => n56, Y => n221);
   U369 : AOI22X1 port map( A => n89, B => regg_213_port, C => regg_197_port, D
                           => n53, Y => n222);
   U371 : AOI22X1 port map( A => n90, B => regg_197_port, C => regg_181_port, D
                           => n53, Y => n223);
   U373 : AOI22X1 port map( A => n90, B => regg_181_port, C => regg_165_port, D
                           => n53, Y => n224);
   U375 : AOI22X1 port map( A => n90, B => regg_165_port, C => regg_149_port, D
                           => n53, Y => n225);
   U377 : AOI22X1 port map( A => n90, B => regg_149_port, C => regg_133_port, D
                           => n53, Y => n226);
   U379 : AOI22X1 port map( A => n90, B => regg_133_port, C => regg_117_port, D
                           => n53, Y => n227);
   U381 : AOI22X1 port map( A => n91, B => regg_117_port, C => regg_101_port, D
                           => n55, Y => n228);
   U383 : AOI22X1 port map( A => regg_85_port, B => n61, C => n75, D => 
                           regg_101_port, Y => n229);
   U385 : AOI22X1 port map( A => n91, B => regg_85_port, C => regg_69_port, D 
                           => n55, Y => n230);
   U387 : AOI22X1 port map( A => n92, B => regg_69_port, C => regg_53_port, D 
                           => n55, Y => n231);
   U389 : AOI22X1 port map( A => n92, B => regg_53_port, C => regg_37_port, D 
                           => n55, Y => n232);
   U390 : OAI22X1 port map( A => n63, B => n789, C => n788, D => n70, Y => n500
                           );
   U392 : OAI22X1 port map( A => n787, B => n78, C => n62, D => n788, Y => n501
                           );
   U394 : OAI21X1 port map( A => n64, B => n787, C => n236, Y => n502);
   U395 : NAND2X1 port map( A => databus_out(5), B => n65, Y => n236);
   U398 : AOI22X1 port map( A => n93, B => regg_246_port, C => regg_230_port, D
                           => n54, Y => n237);
   U400 : AOI22X1 port map( A => n93, B => regg_230_port, C => regg_214_port, D
                           => n54, Y => n238);
   U402 : AOI22X1 port map( A => n93, B => regg_214_port, C => regg_198_port, D
                           => n54, Y => n239);
   U404 : AOI22X1 port map( A => n93, B => regg_198_port, C => regg_182_port, D
                           => n54, Y => n240);
   U406 : AOI22X1 port map( A => n93, B => regg_182_port, C => regg_166_port, D
                           => n54, Y => n241);
   U408 : AOI22X1 port map( A => n94, B => regg_166_port, C => regg_150_port, D
                           => n54, Y => n242);
   U410 : AOI22X1 port map( A => n94, B => regg_150_port, C => regg_134_port, D
                           => n54, Y => n243);
   U412 : AOI22X1 port map( A => n94, B => regg_134_port, C => regg_118_port, D
                           => n53, Y => n244);
   U414 : AOI22X1 port map( A => n95, B => regg_118_port, C => regg_102_port, D
                           => n53, Y => n245);
   U416 : AOI22X1 port map( A => regg_86_port, B => n61, C => n74, D => 
                           regg_102_port, Y => n246);
   U418 : AOI22X1 port map( A => n95, B => regg_86_port, C => regg_70_port, D 
                           => n53, Y => n247);
   U420 : AOI22X1 port map( A => n95, B => regg_70_port, C => regg_54_port, D 
                           => n52, Y => n248);
   U422 : AOI22X1 port map( A => n96, B => regg_54_port, C => regg_38_port, D 
                           => n52, Y => n249);
   U423 : OAI22X1 port map( A => n63, B => n786, C => n785, D => n70, Y => n516
                           );
   U425 : OAI22X1 port map( A => n784, B => n78, C => n62, D => n785, Y => n517
                           );
   U427 : OAI21X1 port map( A => n64, B => n784, C => n253, Y => n518);
   U428 : NAND2X1 port map( A => databus_out(6), B => n64, Y => n253);
   U431 : AOI22X1 port map( A => n89, B => regg_247_port, C => regg_231_port, D
                           => n51, Y => n254);
   U433 : AOI22X1 port map( A => n133, B => regg_231_port, C => regg_215_port, 
                           D => n51, Y => n255);
   U435 : AOI22X1 port map( A => n117, B => regg_215_port, C => regg_199_port, 
                           D => n51, Y => n256);
   U437 : AOI22X1 port map( A => n117, B => regg_199_port, C => regg_183_port, 
                           D => n51, Y => n257);
   U439 : AOI22X1 port map( A => n117, B => regg_183_port, C => regg_167_port, 
                           D => n50, Y => n258);
   U441 : AOI22X1 port map( A => n117, B => regg_167_port, C => regg_151_port, 
                           D => n50, Y => n259);
   U443 : AOI22X1 port map( A => n117, B => regg_151_port, C => regg_135_port, 
                           D => n50, Y => n260);
   U445 : AOI22X1 port map( A => n116, B => regg_135_port, C => regg_119_port, 
                           D => n50, Y => n261);
   U447 : AOI22X1 port map( A => n116, B => regg_119_port, C => regg_103_port, 
                           D => n50, Y => n262);
   U449 : AOI22X1 port map( A => regg_87_port, B => n61, C => n76, D => 
                           regg_103_port, Y => n263);
   U451 : AOI22X1 port map( A => n116, B => regg_87_port, C => regg_71_port, D 
                           => n49, Y => n264);
   U453 : AOI22X1 port map( A => n116, B => regg_71_port, C => regg_55_port, D 
                           => n49, Y => n265);
   U455 : AOI22X1 port map( A => n116, B => regg_55_port, C => regg_39_port, D 
                           => n49, Y => n266);
   U456 : OAI22X1 port map( A => n62, B => n783, C => n782, D => n71, Y => n532
                           );
   U458 : OAI22X1 port map( A => n781, B => n78, C => n62, D => n782, Y => n533
                           );
   U460 : OAI21X1 port map( A => n65, B => n781, C => n270, Y => n534);
   U461 : NAND2X1 port map( A => databus_out(7), B => n65, Y => n270);
   U464 : AOI22X1 port map( A => n115, B => regg_248_port, C => regg_232_port, 
                           D => n48, Y => n271);
   U466 : AOI22X1 port map( A => n115, B => regg_232_port, C => regg_216_port, 
                           D => n48, Y => n272);
   U468 : AOI22X1 port map( A => n115, B => regg_216_port, C => regg_200_port, 
                           D => n48, Y => n273);
   U470 : AOI22X1 port map( A => n115, B => regg_200_port, C => regg_184_port, 
                           D => n47, Y => n274);
   U472 : AOI22X1 port map( A => n115, B => regg_184_port, C => regg_168_port, 
                           D => n47, Y => n275);
   U474 : AOI22X1 port map( A => n114, B => regg_168_port, C => regg_152_port, 
                           D => n47, Y => n276);
   U476 : AOI22X1 port map( A => n114, B => regg_152_port, C => regg_136_port, 
                           D => n46, Y => n277);
   U478 : AOI22X1 port map( A => n114, B => regg_136_port, C => regg_120_port, 
                           D => n46, Y => n278);
   U480 : AOI22X1 port map( A => n114, B => regg_120_port, C => regg_104_port, 
                           D => n46, Y => n279);
   U482 : AOI22X1 port map( A => regg_88_port, B => n60, C => n75, D => 
                           regg_104_port, Y => n280);
   U484 : AOI22X1 port map( A => n114, B => regg_88_port, C => regg_72_port, D 
                           => n57, Y => n281);
   U486 : AOI22X1 port map( A => n113, B => regg_72_port, C => regg_56_port, D 
                           => n57, Y => n282);
   U488 : AOI22X1 port map( A => n113, B => regg_56_port, C => regg_40_port, D 
                           => n57, Y => n283);
   U489 : OAI22X1 port map( A => n64, B => n780, C => n779, D => n72, Y => n548
                           );
   U491 : OAI22X1 port map( A => n778, B => n79, C => n62, D => n779, Y => n549
                           );
   U493 : OAI21X1 port map( A => n65, B => n778, C => n287, Y => n550);
   U494 : NAND2X1 port map( A => databus_out(8), B => n65, Y => n287);
   U497 : AOI22X1 port map( A => n113, B => regg_249_port, C => regg_233_port, 
                           D => n58, Y => n288);
   U499 : AOI22X1 port map( A => n113, B => regg_233_port, C => regg_217_port, 
                           D => n60, Y => n289);
   U501 : AOI22X1 port map( A => n113, B => regg_217_port, C => regg_201_port, 
                           D => n58, Y => n290);
   U503 : AOI22X1 port map( A => n112, B => regg_201_port, C => regg_185_port, 
                           D => n58, Y => n291);
   U505 : AOI22X1 port map( A => n112, B => regg_185_port, C => regg_169_port, 
                           D => n58, Y => n292);
   U507 : AOI22X1 port map( A => n112, B => regg_169_port, C => regg_153_port, 
                           D => n58, Y => n293);
   U509 : AOI22X1 port map( A => n112, B => regg_153_port, C => regg_137_port, 
                           D => n59, Y => n294);
   U511 : AOI22X1 port map( A => n112, B => regg_137_port, C => regg_121_port, 
                           D => n59, Y => n295);
   U513 : AOI22X1 port map( A => n111, B => regg_121_port, C => regg_105_port, 
                           D => n58, Y => n296);
   U515 : AOI22X1 port map( A => regg_89_port, B => n61, C => n76, D => 
                           regg_105_port, Y => n297);
   U517 : AOI22X1 port map( A => n111, B => regg_89_port, C => regg_73_port, D 
                           => n59, Y => n298);
   U519 : AOI22X1 port map( A => n111, B => regg_73_port, C => regg_57_port, D 
                           => n59, Y => n299);
   U521 : AOI22X1 port map( A => n111, B => regg_57_port, C => regg_41_port, D 
                           => n59, Y => n300);
   U522 : OAI22X1 port map( A => n64, B => n777, C => n776, D => n72, Y => n564
                           );
   U524 : OAI22X1 port map( A => n775, B => n78, C => n62, D => n776, Y => n565
                           );
   U526 : OAI21X1 port map( A => n65, B => n775, C => n304, Y => n566);
   U527 : NAND2X1 port map( A => databus_out(9), B => n62, Y => n304);
   U530 : AOI22X1 port map( A => n111, B => regg_250_port, C => regg_234_port, 
                           D => n57, Y => n305);
   U532 : AOI22X1 port map( A => n110, B => regg_234_port, C => regg_218_port, 
                           D => n57, Y => n306);
   U534 : AOI22X1 port map( A => n110, B => regg_218_port, C => regg_202_port, 
                           D => n57, Y => n307);
   U536 : AOI22X1 port map( A => n110, B => regg_202_port, C => regg_186_port, 
                           D => n56, Y => n308);
   U538 : AOI22X1 port map( A => n110, B => regg_186_port, C => regg_170_port, 
                           D => n56, Y => n309);
   U540 : AOI22X1 port map( A => n110, B => regg_170_port, C => regg_154_port, 
                           D => n56, Y => n310);
   U542 : AOI22X1 port map( A => n109, B => regg_154_port, C => regg_138_port, 
                           D => n56, Y => n311);
   U544 : AOI22X1 port map( A => n109, B => regg_138_port, C => regg_122_port, 
                           D => n56, Y => n312);
   U546 : AOI22X1 port map( A => n109, B => regg_122_port, C => regg_106_port, 
                           D => n56, Y => n313);
   U548 : AOI22X1 port map( A => regg_90_port, B => n61, C => n75, D => 
                           regg_106_port, Y => n314);
   U550 : AOI22X1 port map( A => n109, B => regg_90_port, C => regg_74_port, D 
                           => n55, Y => n315);
   U552 : AOI22X1 port map( A => n109, B => regg_74_port, C => regg_58_port, D 
                           => n55, Y => n316);
   U554 : AOI22X1 port map( A => n108, B => regg_58_port, C => regg_42_port, D 
                           => n55, Y => n317);
   U555 : OAI22X1 port map( A => n63, B => n774, C => n773, D => n72, Y => n580
                           );
   U557 : OAI22X1 port map( A => n63, B => n773, C => n772, D => n74, Y => n581
                           );
   U559 : OAI21X1 port map( A => n64, B => n772, C => n321, Y => n582);
   U560 : NAND2X1 port map( A => databus_out(10), B => n61, Y => n321);
   U563 : AOI22X1 port map( A => n108, B => regg_251_port, C => regg_235_port, 
                           D => n54, Y => n322);
   U565 : AOI22X1 port map( A => n108, B => regg_235_port, C => regg_219_port, 
                           D => n54, Y => n323);
   U567 : AOI22X1 port map( A => n108, B => regg_219_port, C => regg_203_port, 
                           D => n54, Y => n324);
   U569 : AOI22X1 port map( A => n108, B => regg_203_port, C => regg_187_port, 
                           D => n54, Y => n325);
   U571 : AOI22X1 port map( A => n107, B => regg_187_port, C => regg_171_port, 
                           D => n53, Y => n326);
   U573 : AOI22X1 port map( A => n107, B => regg_171_port, C => regg_155_port, 
                           D => n53, Y => n327);
   U575 : AOI22X1 port map( A => n107, B => regg_155_port, C => regg_139_port, 
                           D => n52, Y => n328);
   U577 : AOI22X1 port map( A => n107, B => regg_139_port, C => regg_123_port, 
                           D => n52, Y => n329);
   U579 : AOI22X1 port map( A => n106, B => regg_123_port, C => regg_107_port, 
                           D => n51, Y => n330);
   U581 : AOI22X1 port map( A => regg_91_port, B => n61, C => n77, D => 
                           regg_107_port, Y => n331);
   U583 : AOI22X1 port map( A => n106, B => regg_91_port, C => regg_75_port, D 
                           => n51, Y => n332);
   U585 : AOI22X1 port map( A => n106, B => regg_75_port, C => regg_59_port, D 
                           => n50, Y => n333);
   U587 : AOI22X1 port map( A => n106, B => regg_59_port, C => regg_43_port, D 
                           => n50, Y => n334);
   U588 : OAI22X1 port map( A => n63, B => n771, C => n770, D => n74, Y => n596
                           );
   U590 : OAI22X1 port map( A => n63, B => n770, C => n769, D => n73, Y => n597
                           );
   U592 : OAI21X1 port map( A => n64, B => n769, C => n338, Y => n598);
   U593 : NAND2X1 port map( A => databus_out(11), B => n63, Y => n338);
   U596 : AOI22X1 port map( A => n106, B => regg_252_port, C => regg_236_port, 
                           D => n48, Y => n339);
   U598 : AOI22X1 port map( A => n105, B => regg_236_port, C => regg_220_port, 
                           D => n47, Y => n340);
   U600 : AOI22X1 port map( A => n105, B => regg_220_port, C => regg_204_port, 
                           D => n47, Y => n341);
   U602 : AOI22X1 port map( A => n105, B => regg_204_port, C => regg_188_port, 
                           D => n46, Y => n342);
   U604 : AOI22X1 port map( A => n105, B => regg_188_port, C => regg_172_port, 
                           D => n46, Y => n343);
   U606 : AOI22X1 port map( A => n105, B => regg_172_port, C => regg_156_port, 
                           D => n60, Y => n344);
   U608 : AOI22X1 port map( A => n104, B => regg_156_port, C => regg_140_port, 
                           D => n60, Y => n345);
   U610 : AOI22X1 port map( A => n104, B => regg_140_port, C => regg_124_port, 
                           D => n60, Y => n346);
   U612 : AOI22X1 port map( A => n104, B => regg_124_port, C => regg_108_port, 
                           D => n60, Y => n347);
   U614 : AOI22X1 port map( A => regg_92_port, B => n61, C => n77, D => 
                           regg_108_port, Y => n348);
   U616 : AOI22X1 port map( A => n104, B => regg_92_port, C => regg_76_port, D 
                           => n60, Y => n349);
   U618 : AOI22X1 port map( A => n104, B => regg_76_port, C => regg_60_port, D 
                           => n59, Y => n350);
   U620 : AOI22X1 port map( A => n103, B => regg_60_port, C => regg_44_port, D 
                           => n59, Y => n351);
   U621 : OAI22X1 port map( A => n63, B => n768, C => n767, D => n74, Y => n612
                           );
   U623 : OAI22X1 port map( A => n63, B => n767, C => n766, D => n71, Y => n613
                           );
   U625 : OAI21X1 port map( A => n64, B => n766, C => n355, Y => n614);
   U626 : NAND2X1 port map( A => databus_out(12), B => n62, Y => n355);
   U629 : AOI22X1 port map( A => n103, B => regg_253_port, C => regg_237_port, 
                           D => n57, Y => n356);
   U631 : AOI22X1 port map( A => n103, B => regg_237_port, C => regg_221_port, 
                           D => n57, Y => n357);
   U633 : AOI22X1 port map( A => n103, B => regg_221_port, C => regg_205_port, 
                           D => n56, Y => n358);
   U635 : AOI22X1 port map( A => n103, B => regg_205_port, C => regg_189_port, 
                           D => n56, Y => n359);
   U637 : AOI22X1 port map( A => n102, B => regg_189_port, C => regg_173_port, 
                           D => n56, Y => n360);
   U639 : AOI22X1 port map( A => n102, B => regg_173_port, C => regg_157_port, 
                           D => n55, Y => n361);
   U641 : AOI22X1 port map( A => n102, B => regg_157_port, C => regg_141_port, 
                           D => n55, Y => n362);
   U643 : AOI22X1 port map( A => n102, B => regg_141_port, C => regg_125_port, 
                           D => n55, Y => n363);
   U645 : AOI22X1 port map( A => n102, B => regg_125_port, C => regg_109_port, 
                           D => n54, Y => n364);
   U647 : AOI22X1 port map( A => regg_93_port, B => n61, C => n77, D => 
                           regg_109_port, Y => n365);
   U649 : AOI22X1 port map( A => n101, B => regg_93_port, C => regg_77_port, D 
                           => n53, Y => n366);
   U651 : AOI22X1 port map( A => n101, B => regg_77_port, C => regg_61_port, D 
                           => n53, Y => n367);
   U653 : AOI22X1 port map( A => n101, B => regg_61_port, C => regg_45_port, D 
                           => n52, Y => n368);
   U654 : OAI22X1 port map( A => n64, B => n765, C => n764, D => n72, Y => n628
                           );
   U656 : OAI22X1 port map( A => n63, B => n764, C => n763, D => n71, Y => n629
                           );
   U658 : OAI21X1 port map( A => n65, B => n763, C => n372, Y => n630);
   U659 : NAND2X1 port map( A => databus_out(13), B => n65, Y => n372);
   U662 : AOI22X1 port map( A => n101, B => regg_254_port, C => regg_238_port, 
                           D => n48, Y => n373);
   U664 : AOI22X1 port map( A => n101, B => regg_238_port, C => regg_222_port, 
                           D => n47, Y => n374);
   U666 : AOI22X1 port map( A => n100, B => regg_222_port, C => regg_206_port, 
                           D => n46, Y => n375);
   U668 : AOI22X1 port map( A => n100, B => regg_206_port, C => regg_190_port, 
                           D => n60, Y => n376);
   U670 : AOI22X1 port map( A => n100, B => regg_190_port, C => regg_174_port, 
                           D => n60, Y => n377);
   U672 : AOI22X1 port map( A => n100, B => regg_174_port, C => regg_158_port, 
                           D => n60, Y => n378);
   U674 : AOI22X1 port map( A => n100, B => regg_158_port, C => regg_142_port, 
                           D => n59, Y => n379);
   U676 : AOI22X1 port map( A => n99, B => regg_142_port, C => regg_126_port, D
                           => n59, Y => n380);
   U678 : AOI22X1 port map( A => n99, B => regg_126_port, C => regg_110_port, D
                           => n58, Y => n381);
   U680 : AOI22X1 port map( A => regg_94_port, B => n61, C => n76, D => 
                           regg_110_port, Y => n382);
   U682 : AOI22X1 port map( A => n99, B => regg_94_port, C => regg_78_port, D 
                           => n56, Y => n383);
   U684 : AOI22X1 port map( A => n99, B => regg_78_port, C => regg_62_port, D 
                           => n55, Y => n384);
   U686 : AOI22X1 port map( A => n99, B => regg_62_port, C => regg_46_port, D 
                           => n55, Y => n385);
   U687 : OAI22X1 port map( A => n63, B => n762, C => n761, D => n72, Y => n644
                           );
   U689 : OAI22X1 port map( A => n63, B => n761, C => n760, D => n71, Y => n645
                           );
   U691 : OAI21X1 port map( A => n65, B => n760, C => n389, Y => n646);
   U692 : NAND2X1 port map( A => databus_out(14), B => n65, Y => n389);
   U695 : AOI22X1 port map( A => n98, B => regg_255_port, C => regg_239_port, D
                           => n48, Y => n390);
   U697 : AOI22X1 port map( A => n98, B => regg_239_port, C => regg_223_port, D
                           => n46, Y => n391);
   U699 : AOI22X1 port map( A => n98, B => regg_223_port, C => regg_207_port, D
                           => n50, Y => n392);
   U701 : AOI22X1 port map( A => n98, B => regg_207_port, C => regg_191_port, D
                           => n49, Y => n393);
   U703 : AOI22X1 port map( A => n98, B => regg_191_port, C => regg_175_port, D
                           => n58, Y => n394);
   U705 : AOI22X1 port map( A => n97, B => regg_175_port, C => regg_159_port, D
                           => n49, Y => n395);
   U707 : AOI22X1 port map( A => n97, B => regg_159_port, C => regg_143_port, D
                           => n55, Y => n396);
   U709 : AOI22X1 port map( A => n97, B => regg_143_port, C => regg_127_port, D
                           => n57, Y => n397);
   U711 : AOI22X1 port map( A => n97, B => regg_127_port, C => regg_111_port, D
                           => n60, Y => n398);
   U713 : AOI22X1 port map( A => regg_95_port, B => n61, C => n75, D => 
                           regg_111_port, Y => n399);
   U715 : AOI22X1 port map( A => n97, B => regg_95_port, C => regg_79_port, D 
                           => n51, Y => n400);
   U717 : AOI22X1 port map( A => n107, B => regg_79_port, C => regg_63_port, D 
                           => n54, Y => n401);
   U719 : AOI22X1 port map( A => n96, B => regg_63_port, C => regg_47_port, D 
                           => n52, Y => n402);
   U720 : OAI22X1 port map( A => n64, B => n759, C => n758, D => n70, Y => n660
                           );
   U722 : OAI22X1 port map( A => n62, B => n758, C => n757, D => n70, Y => n661
                           );
   U725 : OAI21X1 port map( A => n65, B => n757, C => n406, Y => n662);
   U726 : NAND2X1 port map( A => databus_out(15), B => n65, Y => n406);
   U2 : INVX1 port map( A => n150, Y => n1);
   U3 : BUFX2 port map( A => n37, Y => n2);
   U4 : BUFX2 port map( A => n17, Y => n37);
   U5 : BUFX4 port map( A => n14, Y => n4);
   U6 : BUFX2 port map( A => n12, Y => n3);
   U7 : BUFX2 port map( A => n10, Y => n38);
   U8 : BUFX4 port map( A => n519, Y => n44);
   U9 : BUFX4 port map( A => n10, Y => n39);
   U10 : BUFX2 port map( A => n14, Y => n16);
   U11 : INVX2 port map( A => n15, Y => n17);
   U12 : BUFX4 port map( A => n12, Y => n9);
   U13 : INVX2 port map( A => n167, Y => n515);
   U14 : INVX4 port map( A => n16, Y => n11);
   U15 : BUFX4 port map( A => n514, Y => n36);
   U16 : INVX2 port map( A => n6, Y => n5);
   U17 : INVX4 port map( A => n36, Y => n6);
   U18 : BUFX2 port map( A => n44, Y => n41);
   U19 : BUFX2 port map( A => n35, Y => n34);
   U20 : INVX8 port map( A => n6, Y => n7);
   U21 : INVX8 port map( A => n6, Y => n8);
   U22 : INVX2 port map( A => n167, Y => n10);
   U23 : BUFX4 port map( A => n515, Y => n19);
   U24 : INVX8 port map( A => n11, Y => n12);
   U25 : INVX1 port map( A => n150, Y => n13);
   U26 : INVX4 port map( A => n150, Y => n514);
   U27 : BUFX2 port map( A => n42, Y => n45);
   U28 : INVX2 port map( A => n15, Y => n14);
   U29 : INVX2 port map( A => n166, Y => n32);
   U30 : NAND2X1 port map( A => row_sel(0), B => row_sel(1), Y => n15);
   U31 : INVX2 port map( A => n68, Y => n53);
   U32 : INVX2 port map( A => n69, Y => n47);
   U33 : INVX2 port map( A => n68, Y => n56);
   U34 : INVX2 port map( A => n69, Y => n48);
   U35 : INVX2 port map( A => n69, Y => n50);
   U36 : INVX2 port map( A => n69, Y => n49);
   U37 : INVX2 port map( A => n68, Y => n55);
   U38 : INVX2 port map( A => n69, Y => n51);
   U39 : INVX2 port map( A => n68, Y => n54);
   U40 : INVX2 port map( A => n68, Y => n52);
   U41 : INVX2 port map( A => n67, Y => n59);
   U42 : INVX2 port map( A => n67, Y => n58);
   U43 : INVX2 port map( A => n67, Y => n57);
   U44 : INVX2 port map( A => n67, Y => n60);
   U45 : INVX2 port map( A => n67, Y => n61);
   U46 : INVX2 port map( A => n66, Y => n62);
   U47 : INVX2 port map( A => n66, Y => n63);
   U48 : INVX2 port map( A => n66, Y => n64);
   U49 : INVX2 port map( A => n66, Y => n65);
   U50 : INVX2 port map( A => n70, Y => n46);
   U51 : BUFX2 port map( A => n135, Y => n69);
   U52 : BUFX2 port map( A => n135, Y => n68);
   U53 : BUFX2 port map( A => n148, Y => n67);
   U54 : BUFX2 port map( A => n148, Y => n66);
   U55 : BUFX2 port map( A => n135, Y => n70);
   U56 : BUFX2 port map( A => n133, Y => n73);
   U57 : BUFX2 port map( A => n133, Y => n72);
   U58 : BUFX2 port map( A => n133, Y => n71);
   U59 : BUFX2 port map( A => n132, Y => n74);
   U60 : BUFX2 port map( A => n131, Y => n77);
   U61 : BUFX2 port map( A => n132, Y => n76);
   U62 : BUFX2 port map( A => n132, Y => n75);
   U63 : BUFX2 port map( A => n131, Y => n78);
   U64 : BUFX2 port map( A => n131, Y => n79);
   U65 : BUFX2 port map( A => n130, Y => n80);
   U66 : BUFX2 port map( A => n130, Y => n81);
   U67 : BUFX2 port map( A => n130, Y => n82);
   U68 : BUFX2 port map( A => n129, Y => n83);
   U69 : BUFX2 port map( A => n129, Y => n84);
   U70 : BUFX2 port map( A => n129, Y => n85);
   U71 : BUFX2 port map( A => n128, Y => n86);
   U72 : BUFX2 port map( A => n128, Y => n87);
   U73 : BUFX2 port map( A => n128, Y => n88);
   U74 : BUFX2 port map( A => n127, Y => n90);
   U75 : BUFX2 port map( A => n127, Y => n91);
   U76 : BUFX2 port map( A => n126, Y => n92);
   U77 : BUFX2 port map( A => n126, Y => n93);
   U78 : BUFX2 port map( A => n126, Y => n94);
   U79 : BUFX2 port map( A => n125, Y => n95);
   U80 : BUFX2 port map( A => n127, Y => n89);
   U81 : BUFX2 port map( A => n118, Y => n117);
   U82 : BUFX2 port map( A => n118, Y => n116);
   U83 : BUFX2 port map( A => n119, Y => n115);
   U84 : BUFX2 port map( A => n119, Y => n114);
   U85 : BUFX2 port map( A => n119, Y => n113);
   U86 : BUFX2 port map( A => n120, Y => n112);
   U87 : BUFX2 port map( A => n120, Y => n111);
   U88 : BUFX2 port map( A => n120, Y => n110);
   U89 : BUFX2 port map( A => n121, Y => n109);
   U90 : BUFX2 port map( A => n121, Y => n108);
   U91 : BUFX2 port map( A => n122, Y => n106);
   U92 : BUFX2 port map( A => n122, Y => n105);
   U93 : BUFX2 port map( A => n122, Y => n104);
   U94 : BUFX2 port map( A => n123, Y => n103);
   U95 : BUFX2 port map( A => n123, Y => n102);
   U96 : BUFX2 port map( A => n123, Y => n101);
   U97 : BUFX2 port map( A => n124, Y => n100);
   U98 : BUFX2 port map( A => n124, Y => n99);
   U99 : BUFX2 port map( A => n124, Y => n98);
   U100 : BUFX2 port map( A => n125, Y => n97);
   U101 : BUFX2 port map( A => n121, Y => n107);
   U102 : BUFX2 port map( A => n125, Y => n96);
   U103 : BUFX2 port map( A => n149, Y => n135);
   U104 : BUFX2 port map( A => n149, Y => n148);
   U105 : BUFX2 port map( A => n149, Y => n118);
   U106 : BUFX2 port map( A => n149, Y => n119);
   U107 : BUFX2 port map( A => n118, Y => n120);
   U108 : BUFX2 port map( A => n149, Y => n130);
   U109 : BUFX2 port map( A => n149, Y => n129);
   U110 : BUFX2 port map( A => n149, Y => n128);
   U111 : BUFX2 port map( A => n149, Y => n126);
   U112 : BUFX2 port map( A => n149, Y => n127);
   U113 : BUFX2 port map( A => n119, Y => n122);
   U114 : BUFX2 port map( A => n123, Y => n131);
   U115 : BUFX2 port map( A => n130, Y => n123);
   U116 : BUFX2 port map( A => n129, Y => n124);
   U117 : BUFX2 port map( A => n122, Y => n132);
   U118 : BUFX2 port map( A => n128, Y => n121);
   U119 : BUFX2 port map( A => n126, Y => n125);
   U120 : BUFX2 port map( A => n120, Y => n133);
   U121 : INVX2 port map( A => strb_matrix, Y => n149);
   U122 : BUFX2 port map( A => n514, Y => n35);
   U123 : BUFX2 port map( A => n39, Y => n18);
   U124 : BUFX2 port map( A => n38, Y => n20);
   U125 : BUFX2 port map( A => n38, Y => n21);
   U126 : BUFX2 port map( A => n40, Y => n22);
   U127 : BUFX2 port map( A => n40, Y => n23);
   U128 : BUFX2 port map( A => n40, Y => n24);
   U129 : BUFX2 port map( A => n39, Y => n25);
   U130 : BUFX2 port map( A => n39, Y => n26);
   U131 : BUFX2 port map( A => n38, Y => n27);
   U132 : BUFX2 port map( A => n38, Y => n28);
   U133 : BUFX2 port map( A => n38, Y => n29);
   U134 : BUFX2 port map( A => n38, Y => n30);
   U135 : BUFX2 port map( A => n38, Y => n31);
   U136 : BUFX2 port map( A => n38, Y => n40);
   U137 : INVX2 port map( A => n166, Y => n519);
   U138 : BUFX2 port map( A => n32, Y => n42);
   U139 : BUFX4 port map( A => n13, Y => n33);
   U140 : BUFX4 port map( A => n519, Y => n43);
   U141 : INVX2 port map( A => row_sel(1), Y => n165);
   U142 : OR2X2 port map( A => row_sel(0), B => n165, Y => n150);
   U143 : AOI22X1 port map( A => regg_0_port, B => n9, C => regg_64_port, D => 
                           n33, Y => n183);
   U144 : NAND2X1 port map( A => n165, B => row_sel(0), Y => n166);
   U145 : OR2X2 port map( A => row_sel(0), B => row_sel(1), Y => n167);
   U146 : AOI22X1 port map( A => regg_128_port, B => n43, C => regg_192_port, D
                           => n20, Y => n182);
   U147 : NAND2X1 port map( A => n183, B => n182, Y => row(0));
   U148 : AOI22X1 port map( A => regg_1_port, B => n2, C => regg_65_port, D => 
                           n8, Y => n199);
   U149 : AOI22X1 port map( A => regg_129_port, B => n43, C => regg_193_port, D
                           => n19, Y => n184);
   U150 : NAND2X1 port map( A => n199, B => n184, Y => row(1));
   U151 : AOI22X1 port map( A => regg_2_port, B => n3, C => regg_66_port, D => 
                           n34, Y => n201);
   U152 : AOI22X1 port map( A => regg_130_port, B => n41, C => regg_194_port, D
                           => n30, Y => n200);
   U153 : NAND2X1 port map( A => n201, B => n200, Y => row(2));
   U154 : AOI22X1 port map( A => regg_3_port, B => n9, C => regg_67_port, D => 
                           n7, Y => n217);
   U155 : AOI22X1 port map( A => regg_131_port, B => n45, C => regg_195_port, D
                           => n21, Y => n216);
   U156 : NAND2X1 port map( A => n217, B => n216, Y => row(3));
   U157 : AOI22X1 port map( A => regg_4_port, B => n2, C => regg_68_port, D => 
                           n33, Y => n233);
   U158 : AOI22X1 port map( A => regg_132_port, B => n43, C => regg_196_port, D
                           => n22, Y => n218);
   U159 : NAND2X1 port map( A => n233, B => n218, Y => row(4));
   U160 : AOI22X1 port map( A => regg_5_port, B => n3, C => regg_69_port, D => 
                           n8, Y => n235);
   U161 : AOI22X1 port map( A => regg_133_port, B => n43, C => regg_197_port, D
                           => n30, Y => n234);
   U162 : NAND2X1 port map( A => n235, B => n234, Y => row(5));
   U163 : AOI22X1 port map( A => regg_6_port, B => n9, C => regg_70_port, D => 
                           n33, Y => n251);
   U164 : AOI22X1 port map( A => regg_134_port, B => n41, C => regg_198_port, D
                           => n23, Y => n250);
   U165 : NAND2X1 port map( A => n251, B => n250, Y => row(6));
   U166 : AOI22X1 port map( A => regg_7_port, B => n9, C => regg_71_port, D => 
                           n7, Y => n267);
   U167 : AOI22X1 port map( A => regg_135_port, B => n45, C => regg_199_port, D
                           => n24, Y => n252);
   U168 : NAND2X1 port map( A => n267, B => n252, Y => row(7));
   U169 : AOI22X1 port map( A => regg_8_port, B => n2, C => regg_72_port, D => 
                           n34, Y => n269);
   U170 : AOI22X1 port map( A => regg_136_port, B => n43, C => regg_200_port, D
                           => n30, Y => n268);
   U171 : NAND2X1 port map( A => n269, B => n268, Y => row(8));
   U172 : AOI22X1 port map( A => regg_9_port, B => n9, C => regg_73_port, D => 
                           n33, Y => n285);
   U173 : AOI22X1 port map( A => regg_137_port, B => n41, C => regg_201_port, D
                           => n30, Y => n284);
   U174 : NAND2X1 port map( A => n285, B => n284, Y => row(9));
   U175 : AOI22X1 port map( A => regg_10_port, B => n3, C => regg_74_port, D =>
                           n8, Y => n301);
   U176 : AOI22X1 port map( A => regg_138_port, B => n43, C => regg_202_port, D
                           => n30, Y => n286);
   U177 : NAND2X1 port map( A => n301, B => n286, Y => row(10));
   U178 : AOI22X1 port map( A => regg_11_port, B => n9, C => regg_75_port, D =>
                           n7, Y => n303);
   U179 : AOI22X1 port map( A => regg_139_port, B => n43, C => regg_203_port, D
                           => n25, Y => n302);
   U180 : NAND2X1 port map( A => n303, B => n302, Y => row(11));
   U181 : AOI22X1 port map( A => regg_12_port, B => n2, C => regg_76_port, D =>
                           n33, Y => n319);
   U182 : AOI22X1 port map( A => regg_140_port, B => n45, C => regg_204_port, D
                           => n26, Y => n318);
   U183 : NAND2X1 port map( A => n319, B => n318, Y => row(12));
   U184 : AOI22X1 port map( A => regg_13_port, B => n3, C => regg_77_port, D =>
                           n8, Y => n335);
   U185 : AOI22X1 port map( A => regg_141_port, B => n43, C => regg_205_port, D
                           => n30, Y => n320);
   U186 : NAND2X1 port map( A => n335, B => n320, Y => row(13));
   U187 : AOI22X1 port map( A => regg_14_port, B => n3, C => regg_78_port, D =>
                           n34, Y => n337);
   U188 : AOI22X1 port map( A => regg_142_port, B => n41, C => regg_206_port, D
                           => n30, Y => n336);
   U189 : NAND2X1 port map( A => n337, B => n336, Y => row(14));
   U190 : AOI22X1 port map( A => regg_15_port, B => n3, C => regg_79_port, D =>
                           n7, Y => n353);
   U191 : AOI22X1 port map( A => regg_143_port, B => n45, C => regg_207_port, D
                           => n30, Y => n352);
   U192 : NAND2X1 port map( A => n353, B => n352, Y => row(15));
   U193 : NAND2X1 port map( A => n1, B => regg_80_port, Y => n370);
   U194 : NAND2X1 port map( A => regg_208_port, B => n10, Y => n369);
   U195 : AOI22X1 port map( A => regg_16_port, B => n17, C => regg_144_port, D 
                           => n519, Y => n354);
   U196 : NAND3X1 port map( A => n354, B => n370, C => n369, Y => row(16));
   U197 : AOI22X1 port map( A => n32, B => regg_145_port, C => regg_17_port, D 
                           => n17, Y => n387);
   U198 : NAND2X1 port map( A => regg_209_port, B => n10, Y => n386);
   U199 : NAND2X1 port map( A => n1, B => regg_81_port, Y => n371);
   U201 : NAND3X1 port map( A => n387, B => n386, C => n371, Y => row(17));
   U203 : AOI22X1 port map( A => regg_18_port, B => n4, C => regg_82_port, D =>
                           n35, Y => n403);
   U205 : AOI22X1 port map( A => regg_146_port, B => n42, C => regg_210_port, D
                           => n19, Y => n388);
   U207 : NAND2X1 port map( A => n403, B => n388, Y => row(18));
   U209 : AOI22X1 port map( A => regg_19_port, B => n37, C => regg_83_port, D 
                           => n33, Y => n405);
   U211 : AOI22X1 port map( A => regg_147_port, B => n44, C => regg_211_port, D
                           => n38, Y => n404);
   U213 : NAND2X1 port map( A => n405, B => n404, Y => row(19));
   U215 : AOI22X1 port map( A => regg_20_port, B => n12, C => regg_84_port, D 
                           => n8, Y => n408);
   U217 : AOI22X1 port map( A => regg_148_port, B => n43, C => regg_212_port, D
                           => n21, Y => n407);
   U219 : NAND2X1 port map( A => n408, B => n407, Y => row(20));
   U221 : AOI22X1 port map( A => regg_21_port, B => n9, C => regg_85_port, D =>
                           n8, Y => n410);
   U223 : AOI22X1 port map( A => regg_149_port, B => n43, C => regg_213_port, D
                           => n23, Y => n409);
   U226 : NAND2X1 port map( A => n410, B => n409, Y => row(21));
   U228 : AOI22X1 port map( A => regg_22_port, B => n12, C => regg_86_port, D 
                           => n7, Y => n412);
   U231 : AOI22X1 port map( A => regg_150_port, B => n45, C => regg_214_port, D
                           => n26, Y => n411);
   U232 : NAND2X1 port map( A => n412, B => n411, Y => row(22));
   U234 : AOI22X1 port map( A => regg_23_port, B => n9, C => regg_87_port, D =>
                           n8, Y => n414);
   U236 : AOI22X1 port map( A => regg_151_port, B => n41, C => regg_215_port, D
                           => n25, Y => n413);
   U238 : NAND2X1 port map( A => n414, B => n413, Y => row(23));
   U240 : AOI22X1 port map( A => regg_24_port, B => n37, C => regg_88_port, D 
                           => n34, Y => n416);
   U242 : AOI22X1 port map( A => regg_152_port, B => n43, C => regg_216_port, D
                           => n27, Y => n415);
   U244 : NAND2X1 port map( A => n416, B => n415, Y => row(24));
   U246 : AOI22X1 port map( A => regg_25_port, B => n9, C => regg_89_port, D =>
                           n8, Y => n418);
   U248 : AOI22X1 port map( A => regg_153_port, B => n43, C => regg_217_port, D
                           => n29, Y => n417);
   U250 : NAND2X1 port map( A => n418, B => n417, Y => row(25));
   U252 : AOI22X1 port map( A => regg_26_port, B => n37, C => regg_90_port, D 
                           => n7, Y => n423);
   U254 : AOI22X1 port map( A => regg_154_port, B => n43, C => regg_218_port, D
                           => n31, Y => n419);
   U256 : NAND2X1 port map( A => n423, B => n419, Y => row(26));
   U259 : AOI22X1 port map( A => regg_27_port, B => n9, C => regg_91_port, D =>
                           n33, Y => n425);
   U261 : AOI22X1 port map( A => regg_155_port, B => n41, C => regg_219_port, D
                           => n31, Y => n424);
   U264 : NAND2X1 port map( A => n425, B => n424, Y => row(27));
   U265 : AOI22X1 port map( A => regg_28_port, B => n3, C => regg_92_port, D =>
                           n7, Y => n427);
   U267 : AOI22X1 port map( A => regg_156_port, B => n43, C => regg_220_port, D
                           => n31, Y => n426);
   U269 : NAND2X1 port map( A => n427, B => n426, Y => row(28));
   U271 : AOI22X1 port map( A => regg_29_port, B => n9, C => regg_93_port, D =>
                           n8, Y => n429);
   U273 : AOI22X1 port map( A => regg_157_port, B => n43, C => regg_221_port, D
                           => n30, Y => n428);
   U275 : NAND2X1 port map( A => n429, B => n428, Y => row(29));
   U277 : AOI22X1 port map( A => regg_30_port, B => n9, C => regg_94_port, D =>
                           n7, Y => n431);
   U279 : AOI22X1 port map( A => regg_158_port, B => n43, C => regg_222_port, D
                           => n30, Y => n430);
   U281 : NAND2X1 port map( A => n431, B => n430, Y => row(30));
   U283 : AOI22X1 port map( A => regg_31_port, B => n3, C => regg_95_port, D =>
                           n8, Y => n433);
   U285 : AOI22X1 port map( A => regg_159_port, B => n41, C => regg_223_port, D
                           => n18, Y => n432);
   U287 : NAND2X1 port map( A => n433, B => n432, Y => row(31));
   U289 : NAND2X1 port map( A => n514, B => regg_96_port, Y => n439);
   U292 : NAND2X1 port map( A => regg_224_port, B => n10, Y => n435);
   U294 : AOI22X1 port map( A => regg_32_port, B => n17, C => regg_160_port, D 
                           => n519, Y => n434);
   U297 : NAND3X1 port map( A => n439, B => n434, C => n435, Y => row(32));
   U298 : NAND2X1 port map( A => regg_97_port, B => n13, Y => n442);
   U300 : NAND2X1 port map( A => regg_225_port, B => n10, Y => n441);
   U302 : AOI22X1 port map( A => regg_33_port, B => n17, C => regg_161_port, D 
                           => n519, Y => n440);
   U304 : NAND3X1 port map( A => n442, B => n441, C => n440, Y => row(33));
   U306 : AOI22X1 port map( A => regg_34_port, B => n16, C => regg_98_port, D 
                           => n35, Y => n444);
   U308 : AOI22X1 port map( A => regg_162_port, B => n42, C => regg_226_port, D
                           => n39, Y => n443);
   U310 : NAND2X1 port map( A => n444, B => n443, Y => row(34));
   U312 : AOI22X1 port map( A => regg_35_port, B => n12, C => regg_99_port, D 
                           => n7, Y => n446);
   U314 : AOI22X1 port map( A => regg_163_port, B => n44, C => regg_227_port, D
                           => n18, Y => n445);
   U316 : NAND2X1 port map( A => n446, B => n445, Y => row(35));
   U318 : AOI22X1 port map( A => regg_36_port, B => n12, C => regg_100_port, D 
                           => n34, Y => n448);
   U320 : AOI22X1 port map( A => regg_164_port, B => n41, C => regg_228_port, D
                           => n22, Y => n447);
   U322 : NAND2X1 port map( A => n448, B => n447, Y => row(36));
   U325 : AOI22X1 port map( A => regg_37_port, B => n12, C => regg_101_port, D 
                           => n33, Y => n450);
   U327 : AOI22X1 port map( A => regg_165_port, B => n43, C => regg_229_port, D
                           => n24, Y => n449);
   U330 : NAND2X1 port map( A => n450, B => n449, Y => row(37));
   U331 : AOI22X1 port map( A => regg_38_port, B => n37, C => regg_102_port, D 
                           => n34, Y => n455);
   U333 : AOI22X1 port map( A => regg_166_port, B => n43, C => regg_230_port, D
                           => n26, Y => n451);
   U335 : NAND2X1 port map( A => n455, B => n451, Y => row(38));
   U337 : AOI22X1 port map( A => regg_39_port, B => n12, C => regg_103_port, D 
                           => n7, Y => n457);
   U339 : AOI22X1 port map( A => regg_167_port, B => n45, C => regg_231_port, D
                           => n28, Y => n456);
   U341 : NAND2X1 port map( A => n457, B => n456, Y => row(39));
   U343 : AOI22X1 port map( A => regg_40_port, B => n12, C => regg_104_port, D 
                           => n8, Y => n459);
   U345 : AOI22X1 port map( A => regg_168_port, B => n41, C => regg_232_port, D
                           => n27, Y => n458);
   U347 : NAND2X1 port map( A => n459, B => n458, Y => row(40));
   U349 : AOI22X1 port map( A => regg_41_port, B => n12, C => regg_105_port, D 
                           => n33, Y => n461);
   U351 : AOI22X1 port map( A => regg_169_port, B => n43, C => regg_233_port, D
                           => n29, Y => n460);
   U353 : NAND2X1 port map( A => n461, B => n460, Y => row(41));
   U355 : AOI22X1 port map( A => regg_42_port, B => n12, C => regg_106_port, D 
                           => n34, Y => n463);
   U358 : AOI22X1 port map( A => regg_170_port, B => n45, C => regg_234_port, D
                           => n27, Y => n462);
   U360 : NAND2X1 port map( A => n463, B => n462, Y => row(42));
   U363 : AOI22X1 port map( A => regg_43_port, B => n3, C => regg_107_port, D 
                           => n8, Y => n465);
   U364 : AOI22X1 port map( A => regg_171_port, B => n43, C => regg_235_port, D
                           => n29, Y => n464);
   U366 : NAND2X1 port map( A => n465, B => n464, Y => row(43));
   U368 : AOI22X1 port map( A => regg_44_port, B => n2, C => regg_108_port, D 
                           => n33, Y => n467);
   U370 : AOI22X1 port map( A => regg_172_port, B => n43, C => regg_236_port, D
                           => n31, Y => n466);
   U372 : NAND2X1 port map( A => n467, B => n466, Y => row(44));
   U374 : AOI22X1 port map( A => regg_45_port, B => n3, C => regg_109_port, D 
                           => n8, Y => n472);
   U376 : AOI22X1 port map( A => regg_173_port, B => n41, C => regg_237_port, D
                           => n30, Y => n471);
   U378 : NAND2X1 port map( A => n472, B => n471, Y => row(45));
   U380 : AOI22X1 port map( A => regg_46_port, B => n2, C => regg_110_port, D 
                           => n34, Y => n474);
   U382 : AOI22X1 port map( A => regg_174_port, B => n43, C => regg_238_port, D
                           => n30, Y => n473);
   U384 : NAND2X1 port map( A => n474, B => n473, Y => row(46));
   U386 : AOI22X1 port map( A => regg_47_port, B => n3, C => regg_111_port, D 
                           => n7, Y => n476);
   U388 : AOI22X1 port map( A => regg_175_port, B => n45, C => regg_239_port, D
                           => n30, Y => n475);
   U391 : NAND2X1 port map( A => n476, B => n475, Y => row(47));
   U393 : AOI22X1 port map( A => regg_48_port, B => n14, C => regg_112_port, D 
                           => n514, Y => n478);
   U396 : AOI22X1 port map( A => regg_176_port, B => n32, C => regg_240_port, D
                           => n515, Y => n477);
   U397 : NAND2X1 port map( A => n478, B => n477, Y => row(48));
   U399 : NAND2X1 port map( A => regg_113_port, B => n514, Y => n481);
   U401 : NAND2X1 port map( A => regg_241_port, B => n515, Y => n480);
   U403 : AOI22X1 port map( A => regg_49_port, B => n14, C => n32, D => 
                           regg_177_port, Y => n479);
   U405 : NAND3X1 port map( A => n480, B => n481, C => n479, Y => row(49));
   U407 : AOI22X1 port map( A => n4, B => regg_50_port, C => regg_114_port, D 
                           => n36, Y => n483);
   U409 : AOI22X1 port map( A => n519, B => regg_178_port, C => regg_242_port, 
                           D => n19, Y => n482);
   U411 : NAND2X1 port map( A => n483, B => n482, Y => row(50));
   U413 : AOI22X1 port map( A => regg_51_port, B => n37, C => regg_115_port, D 
                           => n5, Y => n488);
   U415 : AOI22X1 port map( A => regg_179_port, B => n44, C => regg_243_port, D
                           => n38, Y => n487);
   U417 : NAND2X1 port map( A => n488, B => n487, Y => row(51));
   U419 : AOI22X1 port map( A => regg_52_port, B => n12, C => regg_116_port, D 
                           => n33, Y => n490);
   U421 : AOI22X1 port map( A => regg_180_port, B => n44, C => regg_244_port, D
                           => n20, Y => n489);
   U424 : NAND2X1 port map( A => n490, B => n489, Y => row(52));
   U426 : AOI22X1 port map( A => regg_53_port, B => n12, C => regg_117_port, D 
                           => n7, Y => n492);
   U429 : AOI22X1 port map( A => regg_181_port, B => n45, C => regg_245_port, D
                           => n26, Y => n491);
   U430 : NAND2X1 port map( A => n492, B => n491, Y => row(53));
   U432 : AOI22X1 port map( A => regg_54_port, B => n9, C => regg_118_port, D 
                           => n33, Y => n494);
   U434 : AOI22X1 port map( A => regg_182_port, B => n41, C => regg_246_port, D
                           => n25, Y => n493);
   U436 : NAND2X1 port map( A => n494, B => n493, Y => row(54));
   U438 : AOI22X1 port map( A => regg_55_port, B => n37, C => regg_119_port, D 
                           => n33, Y => n496);
   U440 : AOI22X1 port map( A => regg_183_port, B => n43, C => regg_247_port, D
                           => n26, Y => n495);
   U442 : NAND2X1 port map( A => n496, B => n495, Y => row(55));
   U444 : AOI22X1 port map( A => regg_56_port, B => n9, C => regg_120_port, D 
                           => n33, Y => n498);
   U446 : AOI22X1 port map( A => regg_184_port, B => n43, C => regg_248_port, D
                           => n28, Y => n497);
   U448 : NAND2X1 port map( A => n498, B => n497, Y => row(56));
   U450 : AOI22X1 port map( A => regg_57_port, B => n37, C => regg_121_port, D 
                           => n7, Y => n503);
   U452 : AOI22X1 port map( A => regg_185_port, B => n45, C => regg_249_port, D
                           => n28, Y => n499);
   U454 : NAND2X1 port map( A => n503, B => n499, Y => row(57));
   U457 : AOI22X1 port map( A => regg_58_port, B => n9, C => regg_122_port, D 
                           => n33, Y => n505);
   U459 : AOI22X1 port map( A => regg_186_port, B => n41, C => regg_250_port, D
                           => n29, Y => n504);
   U462 : NAND2X1 port map( A => n505, B => n504, Y => row(58));
   U463 : AOI22X1 port map( A => regg_59_port, B => n2, C => regg_123_port, D 
                           => n7, Y => n507);
   U465 : AOI22X1 port map( A => regg_187_port, B => n45, C => regg_251_port, D
                           => n28, Y => n506);
   U467 : NAND2X1 port map( A => n507, B => n506, Y => row(59));
   U469 : AOI22X1 port map( A => regg_60_port, B => n9, C => regg_124_port, D 
                           => n33, Y => n509);
   U471 : AOI22X1 port map( A => regg_188_port, B => n45, C => regg_252_port, D
                           => n30, Y => n508);
   U473 : NAND2X1 port map( A => n509, B => n508, Y => row(60));
   U475 : AOI22X1 port map( A => regg_61_port, B => n2, C => regg_125_port, D 
                           => n34, Y => n511);
   U477 : AOI22X1 port map( A => regg_189_port, B => n43, C => regg_253_port, D
                           => n30, Y => n510);
   U479 : NAND2X1 port map( A => n511, B => n510, Y => row(61));
   U481 : AOI22X1 port map( A => regg_62_port, B => n2, C => regg_126_port, D 
                           => n33, Y => n513);
   U483 : AOI22X1 port map( A => regg_190_port, B => n41, C => regg_254_port, D
                           => n30, Y => n512);
   U485 : NAND2X1 port map( A => n513, B => n512, Y => row(62));
   U487 : AOI22X1 port map( A => regg_63_port, B => n9, C => regg_127_port, D 
                           => n33, Y => n521);
   U490 : AOI22X1 port map( A => regg_191_port, B => n45, C => regg_255_port, D
                           => n30, Y => n520);
   U492 : NAND2X1 port map( A => n521, B => n520, Y => row(63));
   U495 : INVX2 port map( A => n134, Y => n522);
   U496 : INVX2 port map( A => n136, Y => n523);
   U498 : INVX2 port map( A => n137, Y => n524);
   U500 : INVX2 port map( A => n138, Y => n525);
   U502 : INVX2 port map( A => n139, Y => n526);
   U504 : INVX2 port map( A => n140, Y => n527);
   U506 : INVX2 port map( A => n141, Y => n528);
   U508 : INVX2 port map( A => n142, Y => n529);
   U510 : INVX2 port map( A => n143, Y => n530);
   U512 : INVX2 port map( A => n144, Y => n531);
   U514 : INVX2 port map( A => n145, Y => n535);
   U516 : INVX2 port map( A => n146, Y => n536);
   U518 : INVX2 port map( A => n147, Y => n537);
   U520 : INVX2 port map( A => n152, Y => n538);
   U523 : INVX2 port map( A => n153, Y => n539);
   U525 : INVX2 port map( A => n154, Y => n540);
   U528 : INVX2 port map( A => n155, Y => n541);
   U529 : INVX2 port map( A => n156, Y => n542);
   U531 : INVX2 port map( A => n157, Y => n543);
   U533 : INVX2 port map( A => n158, Y => n544);
   U535 : INVX2 port map( A => n159, Y => n545);
   U537 : INVX2 port map( A => n160, Y => n546);
   U539 : INVX2 port map( A => n161, Y => n547);
   U541 : INVX2 port map( A => n162, Y => n551);
   U543 : INVX2 port map( A => n163, Y => n552);
   U545 : INVX2 port map( A => n164, Y => n553);
   U547 : INVX2 port map( A => n169, Y => n554);
   U549 : INVX2 port map( A => n170, Y => n555);
   U551 : INVX2 port map( A => n171, Y => n556);
   U553 : INVX2 port map( A => n172, Y => n557);
   U556 : INVX2 port map( A => n173, Y => n558);
   U558 : INVX2 port map( A => n174, Y => n559);
   U561 : INVX2 port map( A => n175, Y => n560);
   U562 : INVX2 port map( A => n176, Y => n561);
   U564 : INVX2 port map( A => n177, Y => n562);
   U566 : INVX2 port map( A => n178, Y => n563);
   U568 : INVX2 port map( A => n179, Y => n567);
   U570 : INVX2 port map( A => n180, Y => n568);
   U572 : INVX2 port map( A => n181, Y => n569);
   U574 : INVX2 port map( A => n186, Y => n570);
   U576 : INVX2 port map( A => n187, Y => n571);
   U578 : INVX2 port map( A => n188, Y => n572);
   U580 : INVX2 port map( A => n189, Y => n573);
   U582 : INVX2 port map( A => n190, Y => n574);
   U584 : INVX2 port map( A => n191, Y => n575);
   U586 : INVX2 port map( A => n192, Y => n576);
   U589 : INVX2 port map( A => n193, Y => n577);
   U591 : INVX2 port map( A => n194, Y => n578);
   U594 : INVX2 port map( A => n195, Y => n579);
   U595 : INVX2 port map( A => n196, Y => n583);
   U597 : INVX2 port map( A => n197, Y => n584);
   U599 : INVX2 port map( A => n198, Y => n585);
   U601 : INVX2 port map( A => n203, Y => n586);
   U603 : INVX2 port map( A => n204, Y => n587);
   U605 : INVX2 port map( A => n205, Y => n588);
   U607 : INVX2 port map( A => n206, Y => n589);
   U609 : INVX2 port map( A => n207, Y => n590);
   U611 : INVX2 port map( A => n208, Y => n591);
   U613 : INVX2 port map( A => n209, Y => n592);
   U615 : INVX2 port map( A => n210, Y => n593);
   U617 : INVX2 port map( A => n211, Y => n594);
   U619 : INVX2 port map( A => n212, Y => n595);
   U622 : INVX2 port map( A => n213, Y => n599);
   U624 : INVX2 port map( A => n214, Y => n600);
   U627 : INVX2 port map( A => n215, Y => n601);
   U628 : INVX2 port map( A => n220, Y => n602);
   U630 : INVX2 port map( A => n221, Y => n603);
   U632 : INVX2 port map( A => n222, Y => n604);
   U634 : INVX2 port map( A => n223, Y => n605);
   U636 : INVX2 port map( A => n224, Y => n606);
   U638 : INVX2 port map( A => n225, Y => n607);
   U640 : INVX2 port map( A => n226, Y => n608);
   U642 : INVX2 port map( A => n227, Y => n609);
   U644 : INVX2 port map( A => n228, Y => n610);
   U646 : INVX2 port map( A => n229, Y => n611);
   U648 : INVX2 port map( A => n230, Y => n615);
   U650 : INVX2 port map( A => n231, Y => n616);
   U652 : INVX2 port map( A => n232, Y => n617);
   U655 : INVX2 port map( A => n237, Y => n618);
   U657 : INVX2 port map( A => n238, Y => n619);
   U660 : INVX2 port map( A => n239, Y => n620);
   U661 : INVX2 port map( A => n240, Y => n621);
   U663 : INVX2 port map( A => n241, Y => n622);
   U665 : INVX2 port map( A => n242, Y => n623);
   U667 : INVX2 port map( A => n243, Y => n624);
   U669 : INVX2 port map( A => n244, Y => n625);
   U671 : INVX2 port map( A => n245, Y => n626);
   U673 : INVX2 port map( A => n246, Y => n627);
   U675 : INVX2 port map( A => n247, Y => n631);
   U677 : INVX2 port map( A => n248, Y => n632);
   U679 : INVX2 port map( A => n249, Y => n633);
   U681 : INVX2 port map( A => n254, Y => n634);
   U683 : INVX2 port map( A => n255, Y => n635);
   U685 : INVX2 port map( A => n256, Y => n636);
   U688 : INVX2 port map( A => n257, Y => n637);
   U690 : INVX2 port map( A => n258, Y => n638);
   U693 : INVX2 port map( A => n259, Y => n639);
   U694 : INVX2 port map( A => n260, Y => n640);
   U696 : INVX2 port map( A => n261, Y => n641);
   U698 : INVX2 port map( A => n262, Y => n642);
   U700 : INVX2 port map( A => n263, Y => n643);
   U702 : INVX2 port map( A => n264, Y => n647);
   U704 : INVX2 port map( A => n265, Y => n648);
   U706 : INVX2 port map( A => n266, Y => n649);
   U708 : INVX2 port map( A => n271, Y => n650);
   U710 : INVX2 port map( A => n272, Y => n651);
   U712 : INVX2 port map( A => n273, Y => n652);
   U714 : INVX2 port map( A => n274, Y => n653);
   U716 : INVX2 port map( A => n275, Y => n654);
   U718 : INVX2 port map( A => n276, Y => n655);
   U721 : INVX2 port map( A => n277, Y => n656);
   U723 : INVX2 port map( A => n278, Y => n657);
   U724 : INVX2 port map( A => n279, Y => n658);
   U727 : INVX2 port map( A => n280, Y => n659);
   U728 : INVX2 port map( A => n281, Y => n663);
   U729 : INVX2 port map( A => n282, Y => n664);
   U730 : INVX2 port map( A => n283, Y => n665);
   U731 : INVX2 port map( A => n288, Y => n666);
   U732 : INVX2 port map( A => n289, Y => n667);
   U733 : INVX2 port map( A => n290, Y => n668);
   U734 : INVX2 port map( A => n291, Y => n669);
   U735 : INVX2 port map( A => n292, Y => n670);
   U736 : INVX2 port map( A => n293, Y => n671);
   U737 : INVX2 port map( A => n294, Y => n672);
   U738 : INVX2 port map( A => n295, Y => n673);
   U739 : INVX2 port map( A => n296, Y => n674);
   U740 : INVX2 port map( A => n297, Y => n675);
   U741 : INVX2 port map( A => n298, Y => n676);
   U742 : INVX2 port map( A => n299, Y => n677);
   U743 : INVX2 port map( A => n300, Y => n678);
   U744 : INVX2 port map( A => n305, Y => n679);
   U745 : INVX2 port map( A => n306, Y => n680);
   U746 : INVX2 port map( A => n307, Y => n681);
   U747 : INVX2 port map( A => n308, Y => n682);
   U748 : INVX2 port map( A => n309, Y => n683);
   U749 : INVX2 port map( A => n310, Y => n684);
   U750 : INVX2 port map( A => n311, Y => n685);
   U751 : INVX2 port map( A => n312, Y => n686);
   U752 : INVX2 port map( A => n313, Y => n687);
   U753 : INVX2 port map( A => n314, Y => n688);
   U754 : INVX2 port map( A => n315, Y => n689);
   U755 : INVX2 port map( A => n316, Y => n690);
   U756 : INVX2 port map( A => n317, Y => n691);
   U757 : INVX2 port map( A => n322, Y => n692);
   U758 : INVX2 port map( A => n323, Y => n693);
   U759 : INVX2 port map( A => n324, Y => n694);
   U760 : INVX2 port map( A => n325, Y => n695);
   U761 : INVX2 port map( A => n326, Y => n696);
   U762 : INVX2 port map( A => n327, Y => n697);
   U763 : INVX2 port map( A => n328, Y => n698);
   U764 : INVX2 port map( A => n329, Y => n699);
   U765 : INVX2 port map( A => n330, Y => n700);
   U766 : INVX2 port map( A => n331, Y => n701);
   U767 : INVX2 port map( A => n332, Y => n702);
   U768 : INVX2 port map( A => n333, Y => n703);
   U769 : INVX2 port map( A => n334, Y => n704);
   U770 : INVX2 port map( A => n339, Y => n705);
   U771 : INVX2 port map( A => n340, Y => n706);
   U772 : INVX2 port map( A => n341, Y => n707);
   U773 : INVX2 port map( A => n342, Y => n708);
   U774 : INVX2 port map( A => n343, Y => n709);
   U775 : INVX2 port map( A => n344, Y => n710);
   U776 : INVX2 port map( A => n345, Y => n711);
   U777 : INVX2 port map( A => n346, Y => n712);
   U778 : INVX2 port map( A => n347, Y => n713);
   U779 : INVX2 port map( A => n348, Y => n714);
   U780 : INVX2 port map( A => n349, Y => n715);
   U781 : INVX2 port map( A => n350, Y => n716);
   U782 : INVX2 port map( A => n351, Y => n717);
   U783 : INVX2 port map( A => n356, Y => n718);
   U784 : INVX2 port map( A => n357, Y => n719);
   U785 : INVX2 port map( A => n358, Y => n720);
   U786 : INVX2 port map( A => n359, Y => n721);
   U787 : INVX2 port map( A => n360, Y => n722);
   U788 : INVX2 port map( A => n361, Y => n723);
   U789 : INVX2 port map( A => n362, Y => n724);
   U790 : INVX2 port map( A => n363, Y => n725);
   U791 : INVX2 port map( A => n364, Y => n726);
   U792 : INVX2 port map( A => n365, Y => n727);
   U793 : INVX2 port map( A => n366, Y => n728);
   U794 : INVX2 port map( A => n367, Y => n729);
   U795 : INVX2 port map( A => n368, Y => n730);
   U796 : INVX2 port map( A => n373, Y => n731);
   U797 : INVX2 port map( A => n374, Y => n732);
   U798 : INVX2 port map( A => n375, Y => n733);
   U799 : INVX2 port map( A => n376, Y => n734);
   U800 : INVX2 port map( A => n377, Y => n735);
   U801 : INVX2 port map( A => n378, Y => n736);
   U802 : INVX2 port map( A => n379, Y => n737);
   U803 : INVX2 port map( A => n380, Y => n738);
   U804 : INVX2 port map( A => n381, Y => n739);
   U805 : INVX2 port map( A => n382, Y => n740);
   U806 : INVX2 port map( A => n383, Y => n741);
   U807 : INVX2 port map( A => n384, Y => n742);
   U808 : INVX2 port map( A => n385, Y => n743);
   U809 : INVX2 port map( A => n390, Y => n744);
   U810 : INVX2 port map( A => n391, Y => n745);
   U811 : INVX2 port map( A => n392, Y => n746);
   U812 : INVX2 port map( A => n393, Y => n747);
   U813 : INVX2 port map( A => n394, Y => n748);
   U814 : INVX2 port map( A => n395, Y => n749);
   U815 : INVX2 port map( A => n396, Y => n750);
   U816 : INVX2 port map( A => n397, Y => n751);
   U817 : INVX2 port map( A => n398, Y => n752);
   U818 : INVX2 port map( A => n399, Y => n753);
   U819 : INVX2 port map( A => n400, Y => n754);
   U820 : INVX2 port map( A => n401, Y => n755);
   U821 : INVX2 port map( A => n402, Y => n756);
   U822 : INVX2 port map( A => regg_15_port, Y => n757);
   U823 : INVX2 port map( A => regg_31_port, Y => n758);
   U824 : INVX2 port map( A => regg_47_port, Y => n759);
   U825 : INVX2 port map( A => regg_14_port, Y => n760);
   U826 : INVX2 port map( A => regg_30_port, Y => n761);
   U827 : INVX2 port map( A => regg_46_port, Y => n762);
   U828 : INVX2 port map( A => regg_13_port, Y => n763);
   U829 : INVX2 port map( A => regg_29_port, Y => n764);
   U830 : INVX2 port map( A => regg_45_port, Y => n765);
   U831 : INVX2 port map( A => regg_12_port, Y => n766);
   U832 : INVX2 port map( A => regg_28_port, Y => n767);
   U833 : INVX2 port map( A => regg_44_port, Y => n768);
   U834 : INVX2 port map( A => regg_11_port, Y => n769);
   U835 : INVX2 port map( A => regg_27_port, Y => n770);
   U836 : INVX2 port map( A => regg_43_port, Y => n771);
   U837 : INVX2 port map( A => regg_10_port, Y => n772);
   U838 : INVX2 port map( A => regg_26_port, Y => n773);
   U839 : INVX2 port map( A => regg_42_port, Y => n774);
   U840 : INVX2 port map( A => regg_9_port, Y => n775);
   U841 : INVX2 port map( A => regg_25_port, Y => n776);
   U842 : INVX2 port map( A => regg_41_port, Y => n777);
   U843 : INVX2 port map( A => regg_8_port, Y => n778);
   U844 : INVX2 port map( A => regg_24_port, Y => n779);
   U845 : INVX2 port map( A => regg_40_port, Y => n780);
   U846 : INVX2 port map( A => regg_7_port, Y => n781);
   U847 : INVX2 port map( A => regg_23_port, Y => n782);
   U848 : INVX2 port map( A => regg_39_port, Y => n783);
   U849 : INVX2 port map( A => regg_6_port, Y => n784);
   U850 : INVX2 port map( A => regg_22_port, Y => n785);
   U851 : INVX2 port map( A => regg_38_port, Y => n786);
   U852 : INVX2 port map( A => regg_5_port, Y => n787);
   U853 : INVX2 port map( A => regg_21_port, Y => n788);
   U854 : INVX2 port map( A => regg_37_port, Y => n789);
   U855 : INVX2 port map( A => regg_4_port, Y => n790);
   U856 : INVX2 port map( A => regg_20_port, Y => n791);
   U857 : INVX2 port map( A => regg_36_port, Y => n792);
   U858 : INVX2 port map( A => regg_3_port, Y => n793);
   U859 : INVX2 port map( A => regg_19_port, Y => n794);
   U860 : INVX2 port map( A => regg_35_port, Y => n795);
   U861 : INVX2 port map( A => regg_2_port, Y => n796);
   U862 : INVX2 port map( A => regg_18_port, Y => n797);
   U863 : INVX2 port map( A => regg_34_port, Y => n798);
   U864 : INVX2 port map( A => regg_1_port, Y => n799);
   U865 : INVX2 port map( A => regg_17_port, Y => n800);
   U866 : INVX2 port map( A => regg_33_port, Y => n801);
   U867 : INVX2 port map( A => regg_0_port, Y => n802);
   U868 : INVX2 port map( A => regg_16_port, Y => n803);
   U869 : INVX2 port map( A => regg_32_port, Y => n804);

end SYN_behavorial;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity screen_buffer is

   port( clk, strb_screen : in std_logic;  screen_cor : in std_logic_vector (7 
         downto 0);  X0, X1, Y0, Y1 : out std_logic_vector (7 downto 0));

end screen_buffer;

architecture SYN_beh of screen_buffer is

   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;
   
   signal X0_7_port, X0_6_port, X0_5_port, X0_4_port, X0_3_port, X0_2_port, 
      X0_1_port, X0_0_port, X1_7_port, X1_6_port, X1_5_port, X1_4_port, 
      X1_3_port, X1_2_port, X1_1_port, X1_0_port, Y0_7_port, Y0_6_port, 
      Y0_5_port, Y0_4_port, Y0_3_port, Y0_2_port, Y0_1_port, Y0_0_port, 
      Y1_7_port, Y1_6_port, Y1_5_port, Y1_4_port, Y1_3_port, Y1_2_port, 
      Y1_1_port, Y1_0_port, n3, n8, n13, n18, n23, n28, n33, n38, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73
      , n1, n2, n4, n5, n6, n7, n9, n10, n11, n12, n14, n15, n16, n17, n19, n20
      , n21, n22, n24, n25, n26, n27, n29, n30, n31, n32, n34, n35, n36, n37, 
      n39, n40, n41, n74, n75 : std_logic;

begin
   X0 <= ( X0_7_port, X0_6_port, X0_5_port, X0_4_port, X0_3_port, X0_2_port, 
      X0_1_port, X0_0_port );
   X1 <= ( X1_7_port, X1_6_port, X1_5_port, X1_4_port, X1_3_port, X1_2_port, 
      X1_1_port, X1_0_port );
   Y0 <= ( Y0_7_port, Y0_6_port, Y0_5_port, Y0_4_port, Y0_3_port, Y0_2_port, 
      Y0_1_port, Y0_0_port );
   Y1 <= ( Y1_7_port, Y1_6_port, Y1_5_port, Y1_4_port, Y1_3_port, Y1_2_port, 
      Y1_1_port, Y1_0_port );
   
   reg1_reg_7_inst : DFFPOSX1 port map( D => n73, CLK => clk, Q => Y1_7_port);
   reg1_reg_15_inst : DFFPOSX1 port map( D => n72, CLK => clk, Q => Y0_7_port);
   reg1_reg_23_inst : DFFPOSX1 port map( D => n71, CLK => clk, Q => X1_7_port);
   reg1_reg_31_inst : DFFPOSX1 port map( D => n70, CLK => clk, Q => X0_7_port);
   reg1_reg_6_inst : DFFPOSX1 port map( D => n69, CLK => clk, Q => Y1_6_port);
   reg1_reg_14_inst : DFFPOSX1 port map( D => n68, CLK => clk, Q => Y0_6_port);
   reg1_reg_22_inst : DFFPOSX1 port map( D => n67, CLK => clk, Q => X1_6_port);
   reg1_reg_30_inst : DFFPOSX1 port map( D => n66, CLK => clk, Q => X0_6_port);
   reg1_reg_5_inst : DFFPOSX1 port map( D => n65, CLK => clk, Q => Y1_5_port);
   reg1_reg_13_inst : DFFPOSX1 port map( D => n64, CLK => clk, Q => Y0_5_port);
   reg1_reg_21_inst : DFFPOSX1 port map( D => n63, CLK => clk, Q => X1_5_port);
   reg1_reg_29_inst : DFFPOSX1 port map( D => n62, CLK => clk, Q => X0_5_port);
   reg1_reg_4_inst : DFFPOSX1 port map( D => n61, CLK => clk, Q => Y1_4_port);
   reg1_reg_12_inst : DFFPOSX1 port map( D => n60, CLK => clk, Q => Y0_4_port);
   reg1_reg_20_inst : DFFPOSX1 port map( D => n59, CLK => clk, Q => X1_4_port);
   reg1_reg_28_inst : DFFPOSX1 port map( D => n58, CLK => clk, Q => X0_4_port);
   reg1_reg_3_inst : DFFPOSX1 port map( D => n57, CLK => clk, Q => Y1_3_port);
   reg1_reg_11_inst : DFFPOSX1 port map( D => n56, CLK => clk, Q => Y0_3_port);
   reg1_reg_19_inst : DFFPOSX1 port map( D => n55, CLK => clk, Q => X1_3_port);
   reg1_reg_27_inst : DFFPOSX1 port map( D => n54, CLK => clk, Q => X0_3_port);
   reg1_reg_2_inst : DFFPOSX1 port map( D => n53, CLK => clk, Q => Y1_2_port);
   reg1_reg_10_inst : DFFPOSX1 port map( D => n52, CLK => clk, Q => Y0_2_port);
   reg1_reg_18_inst : DFFPOSX1 port map( D => n51, CLK => clk, Q => X1_2_port);
   reg1_reg_26_inst : DFFPOSX1 port map( D => n50, CLK => clk, Q => X0_2_port);
   reg1_reg_1_inst : DFFPOSX1 port map( D => n49, CLK => clk, Q => Y1_1_port);
   reg1_reg_9_inst : DFFPOSX1 port map( D => n48, CLK => clk, Q => Y0_1_port);
   reg1_reg_17_inst : DFFPOSX1 port map( D => n47, CLK => clk, Q => X1_1_port);
   reg1_reg_25_inst : DFFPOSX1 port map( D => n46, CLK => clk, Q => X0_1_port);
   reg1_reg_0_inst : DFFPOSX1 port map( D => n45, CLK => clk, Q => Y1_0_port);
   reg1_reg_8_inst : DFFPOSX1 port map( D => n44, CLK => clk, Q => Y0_0_port);
   reg1_reg_16_inst : DFFPOSX1 port map( D => n43, CLK => clk, Q => X1_0_port);
   reg1_reg_24_inst : DFFPOSX1 port map( D => n42, CLK => clk, Q => X0_0_port);
   U2 : OAI21X1 port map( A => n75, B => n1, C => n3, Y => n42);
   U3 : NAND2X1 port map( A => X0_0_port, B => n1, Y => n3);
   U4 : OAI22X1 port map( A => n1, B => n74, C => n2, D => n75, Y => n43);
   U6 : OAI22X1 port map( A => n1, B => n41, C => n2, D => n74, Y => n44);
   U11 : OAI21X1 port map( A => n1, B => n40, C => n8, Y => n46);
   U12 : NAND2X1 port map( A => X0_1_port, B => n1, Y => n8);
   U13 : OAI22X1 port map( A => n1, B => n39, C => n2, D => n40, Y => n47);
   U15 : OAI22X1 port map( A => n1, B => n37, C => n2, D => n39, Y => n48);
   U20 : OAI21X1 port map( A => n1, B => n36, C => n13, Y => n50);
   U21 : NAND2X1 port map( A => X0_2_port, B => n1, Y => n13);
   U22 : OAI22X1 port map( A => n1, B => n35, C => n2, D => n36, Y => n51);
   U24 : OAI22X1 port map( A => n1, B => n34, C => n2, D => n35, Y => n52);
   U29 : OAI21X1 port map( A => n1, B => n32, C => n18, Y => n54);
   U30 : NAND2X1 port map( A => X0_3_port, B => n1, Y => n18);
   U31 : OAI22X1 port map( A => n1, B => n31, C => n2, D => n32, Y => n55);
   U33 : OAI22X1 port map( A => n1, B => n30, C => n2, D => n31, Y => n56);
   U38 : OAI21X1 port map( A => n1, B => n29, C => n23, Y => n58);
   U39 : NAND2X1 port map( A => X0_4_port, B => n1, Y => n23);
   U40 : OAI22X1 port map( A => n1, B => n27, C => n4, D => n29, Y => n59);
   U42 : OAI22X1 port map( A => n1, B => n26, C => n4, D => n27, Y => n60);
   U47 : OAI21X1 port map( A => n1, B => n25, C => n28, Y => n62);
   U48 : NAND2X1 port map( A => X0_5_port, B => n1, Y => n28);
   U49 : OAI22X1 port map( A => n1, B => n24, C => n4, D => n25, Y => n63);
   U51 : OAI22X1 port map( A => n1, B => n22, C => n4, D => n24, Y => n64);
   U56 : OAI21X1 port map( A => n1, B => n21, C => n33, Y => n66);
   U57 : NAND2X1 port map( A => X0_6_port, B => n1, Y => n33);
   U58 : OAI22X1 port map( A => n1, B => n20, C => n4, D => n21, Y => n67);
   U60 : OAI22X1 port map( A => n1, B => n19, C => n4, D => n20, Y => n68);
   U65 : OAI21X1 port map( A => n1, B => n17, C => n38, Y => n70);
   U66 : NAND2X1 port map( A => X0_7_port, B => n1, Y => n38);
   U67 : OAI22X1 port map( A => n1, B => n16, C => n4, D => n17, Y => n71);
   U69 : OAI22X1 port map( A => n1, B => n15, C => n2, D => n16, Y => n72);
   U5 : INVX4 port map( A => strb_screen, Y => n1);
   U7 : MUX2X1 port map( B => n14, A => n15, S => n1, Y => n73);
   U8 : BUFX2 port map( A => strb_screen, Y => n2);
   U9 : BUFX2 port map( A => strb_screen, Y => n4);
   U10 : INVX2 port map( A => Y1_7_port, Y => n15);
   U14 : INVX2 port map( A => Y1_6_port, Y => n19);
   U16 : INVX2 port map( A => Y1_5_port, Y => n22);
   U17 : INVX2 port map( A => Y1_4_port, Y => n26);
   U18 : INVX2 port map( A => Y1_3_port, Y => n30);
   U19 : INVX2 port map( A => Y1_2_port, Y => n34);
   U23 : INVX2 port map( A => Y1_1_port, Y => n37);
   U25 : INVX2 port map( A => Y1_0_port, Y => n41);
   U26 : INVX2 port map( A => screen_cor(0), Y => n5);
   U27 : MUX2X1 port map( B => n41, A => n5, S => n4, Y => n45);
   U28 : INVX2 port map( A => screen_cor(1), Y => n6);
   U32 : MUX2X1 port map( B => n37, A => n6, S => n2, Y => n49);
   U34 : INVX2 port map( A => screen_cor(2), Y => n7);
   U35 : MUX2X1 port map( B => n34, A => n7, S => n4, Y => n53);
   U36 : INVX2 port map( A => screen_cor(3), Y => n9);
   U37 : MUX2X1 port map( B => n30, A => n9, S => n4, Y => n57);
   U41 : INVX2 port map( A => screen_cor(4), Y => n10);
   U43 : MUX2X1 port map( B => n26, A => n10, S => n4, Y => n61);
   U44 : INVX2 port map( A => screen_cor(5), Y => n11);
   U45 : MUX2X1 port map( B => n22, A => n11, S => n2, Y => n65);
   U46 : INVX2 port map( A => screen_cor(6), Y => n12);
   U50 : MUX2X1 port map( B => n19, A => n12, S => n2, Y => n69);
   U52 : INVX2 port map( A => screen_cor(7), Y => n14);
   U53 : INVX2 port map( A => Y0_7_port, Y => n16);
   U54 : INVX2 port map( A => X1_7_port, Y => n17);
   U55 : INVX2 port map( A => Y0_6_port, Y => n20);
   U59 : INVX2 port map( A => X1_6_port, Y => n21);
   U61 : INVX2 port map( A => Y0_5_port, Y => n24);
   U62 : INVX2 port map( A => X1_5_port, Y => n25);
   U63 : INVX2 port map( A => Y0_4_port, Y => n27);
   U64 : INVX2 port map( A => X1_4_port, Y => n29);
   U68 : INVX2 port map( A => Y0_3_port, Y => n31);
   U70 : INVX2 port map( A => X1_3_port, Y => n32);
   U71 : INVX2 port map( A => Y0_2_port, Y => n35);
   U72 : INVX2 port map( A => X1_2_port, Y => n36);
   U73 : INVX2 port map( A => Y0_1_port, Y => n39);
   U74 : INVX2 port map( A => X1_1_port, Y => n40);
   U75 : INVX2 port map( A => Y0_0_port, Y => n74);
   U76 : INVX2 port map( A => X1_0_port, Y => n75);

end SYN_beh;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity Rasterizer is

   port( clk : in std_logic;  X0, X1, Y0, Y1 : in std_logic_vector (7 downto 0)
         ;  init_rast, RST_N : in std_logic;  rast_done, rast_strb : out 
         std_logic;  rast_index : out std_logic_vector (3 downto 0);  rast_addr
         : out std_logic_vector (15 downto 0));

end Rasterizer;

architecture SYN_Mixed of Rasterizer is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AOI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component Rasterizer_DW01_add_3
      port( A, B : in std_logic_vector (8 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (8 downto 0);  CO : out std_logic);
   end component;
   
   component Rasterizer_DW01_sub_6
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  DIFF 
            : out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component Rasterizer_DW01_sub_5
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  DIFF 
            : out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component Rasterizer_DW01_sub_4
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  DIFF 
            : out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component Rasterizer_DW01_sub_3
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  DIFF 
            : out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component Rasterizer_DW01_inc_2
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component Rasterizer_DW01_sub_2
      port( A, B : in std_logic_vector (11 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (11 downto 0);  CO : out std_logic);
   end component;
   
   component Rasterizer_DW01_inc_1
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component Rasterizer_DW01_add_0
      port( A, B : in std_logic_vector (11 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (11 downto 0);  CO : out std_logic);
   end component;
   
   component Rasterizer_DW01_inc_0
      port( A : in std_logic_vector (7 downto 0);  SUM : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI22X1
      port( A, B, C, D : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal rast_index_3_port, rast_index_2_port, rast_index_1_port, 
      rast_index_0_port, rast_addr_11_port, rast_addr_10_port, rast_addr_9_port
      , rast_addr_8_port, rast_addr_7_port, rast_addr_6_port, rast_addr_5_port,
      rast_addr_4_port, rast_addr_3_port, rast_addr_2_port, rast_addr_1_port, 
      rast_addr_0_port, state_3_port, state_2_port, state_1_port, state_0_port,
      dx_8_port, dx_7_port, dx_6_port, dx_5_port, dx_4_port, dx_3_port, 
      dx_2_port, dx_0_port, dy_8_port, dy_7_port, dy_6_port, dy_5_port, 
      dy_4_port, dy_3_port, dy_2_port, dy_1_port, dy_0_port, iX, iY, steep, 
      err_11_port, err_10_port, err_9_port, err_8_port, err_7_port, err_6_port,
      err_5_port, err_4_port, err_3_port, err_2_port, err_1_port, err_0_port, 
      i_7_port, i_6_port, i_5_port, i_4_port, i_3_port, i_2_port, i_1_port, 
      i_0_port, count_3_port, count_2_port, count_1_port, count_0_port, 
      nextstate_3_port, nextstate_2_port, nextstate_1_port, nextstate_0_port, 
      N95, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108,
      N109, N110, N111, N112, N121, N123, N124, N125, N126, N127, N128, N129, 
      N130, N131, N132, N133, N134, N135, N136, N137, N138, N188, N199, N200, 
      N201, N202, N203, N204, N205, N206, N207, N209, N210, N211, N212, N213, 
      N214, N215, N216, N217, N218, N219, N220, N229, N230, N231, N232, N257, 
      N258, N259, N260, N261, N262, N263, N264, N265, N266, N269, N270, N271, 
      N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, 
      N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, 
      N296, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, 
      N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, 
      N329, N330, N331, N332, N333, n3, n4, n13, n14, n16, n17, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95_port, n96, n97_port, 
      n98_port, n99_port, n100_port, n101_port, n102_port, n103_port, n104_port
      , n105_port, n106_port, n107_port, n108_port, n109_port, n110_port, 
      n111_port, n112_port, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121_port, n122, n123_port, n124_port, n125_port, n126_port, n127_port, 
      n128_port, n129_port, n130_port, n131_port, n132_port, n133_port, 
      n134_port, n135_port, n136_port, n137_port, n138_port, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n229_port, n230_port, n231_port
      , n232_port, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257_port, n258_port, n259_port, n260_port, n261_port, 
      n262_port, n263_port, n266_port, n267, n268, n269_port, n270_port, 
      n271_port, n272_port, n273_port, n274_port, n275_port, n276_port, 
      n277_port, n278_port, n279_port, n280_port, n281_port, n282_port, 
      n283_port, n284_port, n285_port, n286_port, n287_port, n288_port, 
      n289_port, n290_port, n291_port, n292_port, n293_port, n294_port, 
      n295_port, n296_port, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306_port, n307_port, n308_port, n309_port, n310_port, n311_port, 
      n312_port, n313_port, n314_port, n315_port, n316_port, n317_port, 
      n318_port, n319_port, n320_port, n321_port, n322_port, n323_port, 
      n324_port, n325_port, n326_port, n327_port, n328_port, n329_port, 
      n330_port, n331_port, n332_port, n333_port, n334, n335, n336, n337, n338,
      n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
      n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, N198, N197, N196, 
      N195, N194, N193, N192, N191, N190, 
      sub_1_root_sub_0_root_sub_184_carry_2_port, 
      sub_1_root_sub_0_root_sub_184_carry_3_port, 
      sub_1_root_sub_0_root_sub_184_carry_4_port, 
      sub_1_root_sub_0_root_sub_184_carry_5_port, 
      sub_1_root_sub_0_root_sub_184_carry_6_port, 
      sub_1_root_sub_0_root_sub_184_carry_7_port, n1, n2, n5, n6, n7, n8, n9, 
      n10, n11, n12, n15, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188_port, n189, n190_port, n191_port, n192_port, n193_port, n194_port, 
      n195_port, n196_port, n197_port, n198_port, n199_port, n200_port, 
      n201_port, n202_port, n203_port, n204_port, n205_port, n206_port, 
      n207_port, n208, n209_port, n210_port, n211_port, n212_port, n213_port, 
      n214_port, n215_port, n216_port, n217_port, n218_port, n219_port, 
      n220_port, n221, n222, n223, n224, n225, n226, n227, n228, n264_port, 
      n265_port, n361, n362, n398, n399, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, 
      rast_done_port, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230 : 
      std_logic;

begin
   rast_done <= rast_done_port;
   rast_index <= ( rast_index_3_port, rast_index_2_port, rast_index_1_port, 
      rast_index_0_port );
   rast_addr <= ( n644, n644, n644, n644, rast_addr_11_port, rast_addr_10_port,
      rast_addr_9_port, rast_addr_8_port, rast_addr_7_port, rast_addr_6_port, 
      rast_addr_5_port, rast_addr_4_port, rast_addr_3_port, rast_addr_2_port, 
      rast_addr_1_port, rast_addr_0_port );
   
   n644 <= '0';
   n3 <= '0';
   n4 <= '0';
   n13 <= '0';
   n14 <= '0';
   n16 <= '0';
   n17 <= '0';
   i_reg_0_inst : DFFSR port map( D => n567, CLK => clk, R => n24, S => n148, Q
                           => i_0_port);
   state_reg_2_inst : DFFSR port map( D => nextstate_2_port, CLK => clk, R => 
                           n21, S => n147, Q => state_2_port);
   dx_reg_0_inst : DFFSR port map( D => n529, CLK => clk, R => n21, S => n146, 
                           Q => dx_0_port);
   dx_reg_1_inst : DFFSR port map( D => n528, CLK => clk, R => n21, S => n145, 
                           Q => N190);
   dx_reg_2_inst : DFFSR port map( D => n527, CLK => clk, R => n21, S => n144, 
                           Q => dx_2_port);
   dx_reg_3_inst : DFFSR port map( D => n526, CLK => clk, R => n21, S => n143, 
                           Q => dx_3_port);
   dx_reg_4_inst : DFFSR port map( D => n525, CLK => clk, R => n21, S => n142, 
                           Q => dx_4_port);
   dx_reg_5_inst : DFFSR port map( D => n524, CLK => clk, R => n21, S => n141, 
                           Q => dx_5_port);
   dx_reg_6_inst : DFFSR port map( D => n523, CLK => clk, R => n21, S => n140, 
                           Q => dx_6_port);
   dx_reg_7_inst : DFFSR port map( D => n522, CLK => clk, R => n21, S => n139, 
                           Q => dx_7_port);
   dx_reg_8_inst : DFFSR port map( D => n521, CLK => clk, R => n21, S => 
                           n138_port, Q => dx_8_port);
   dy_reg_8_inst : DFFSR port map( D => n530, CLK => clk, R => n21, S => 
                           n137_port, Q => dy_8_port);
   dy_reg_7_inst : DFFSR port map( D => n531, CLK => clk, R => n22, S => 
                           n136_port, Q => dy_7_port);
   err_reg_11_inst : DFFSR port map( D => n554, CLK => clk, R => n22, S => 
                           n135_port, Q => err_11_port);
   err_reg_10_inst : DFFSR port map( D => n549, CLK => clk, R => n22, S => 
                           n134_port, Q => err_10_port);
   state_reg_1_inst : DFFSR port map( D => nextstate_1_port, CLK => clk, R => 
                           n22, S => n133_port, Q => state_1_port);
   state_reg_0_inst : DFFSR port map( D => nextstate_0_port, CLK => clk, R => 
                           n22, S => n132_port, Q => state_0_port);
   count_reg_3_inst : DFFSR port map( D => n550, CLK => clk, R => n22, S => 
                           n131_port, Q => count_3_port);
   state_reg_3_inst : DFFSR port map( D => nextstate_3_port, CLK => clk, R => 
                           n22, S => n130_port, Q => state_3_port);
   dy_reg_0_inst : DFFSR port map( D => n538, CLK => clk, R => n22, S => 
                           n129_port, Q => dy_0_port);
   dy_reg_1_inst : DFFSR port map( D => n537, CLK => clk, R => n22, S => 
                           n128_port, Q => dy_1_port);
   dy_reg_2_inst : DFFSR port map( D => n536, CLK => clk, R => n22, S => 
                           n127_port, Q => dy_2_port);
   dy_reg_3_inst : DFFSR port map( D => n535, CLK => clk, R => n22, S => 
                           n126_port, Q => dy_3_port);
   dy_reg_4_inst : DFFSR port map( D => n534, CLK => clk, R => n22, S => 
                           n125_port, Q => dy_4_port);
   dy_reg_5_inst : DFFSR port map( D => n533, CLK => clk, R => n23, S => 
                           n124_port, Q => dy_5_port);
   dy_reg_6_inst : DFFSR port map( D => n532, CLK => clk, R => n23, S => 
                           n123_port, Q => dy_6_port);
   count_reg_0_inst : DFFSR port map( D => n553, CLK => clk, R => n23, S => 
                           n122, Q => count_0_port);
   count_reg_1_inst : DFFSR port map( D => n552, CLK => clk, R => n23, S => 
                           n121_port, Q => count_1_port);
   count_reg_2_inst : DFFSR port map( D => n551, CLK => clk, R => n23, S => 
                           n120, Q => count_2_port);
   iX_reg : DFFSR port map( D => n519, CLK => clk, R => n23, S => n119, Q => iX
                           );
   iY_reg : DFFSR port map( D => n520, CLK => clk, R => n23, S => n118, Q => iY
                           );
   err_reg_9_inst : DFFSR port map( D => n548, CLK => clk, R => n23, S => n117,
                           Q => err_9_port);
   err_reg_8_inst : DFFSR port map( D => n555, CLK => clk, R => n116, S => n27,
                           Q => err_8_port);
   err_reg_7_inst : DFFSR port map( D => n547, CLK => clk, R => n23, S => n115,
                           Q => err_7_port);
   err_reg_6_inst : DFFSR port map( D => n546, CLK => clk, R => n23, S => n114,
                           Q => err_6_port);
   err_reg_5_inst : DFFSR port map( D => n545, CLK => clk, R => n23, S => n113,
                           Q => err_5_port);
   err_reg_4_inst : DFFSR port map( D => n544, CLK => clk, R => n23, S => 
                           n112_port, Q => err_4_port);
   err_reg_3_inst : DFFSR port map( D => n543, CLK => clk, R => n24, S => 
                           n111_port, Q => err_3_port);
   err_reg_2_inst : DFFSR port map( D => n542, CLK => clk, R => n24, S => 
                           n110_port, Q => err_2_port);
   err_reg_1_inst : DFFSR port map( D => n541, CLK => clk, R => n24, S => 
                           n109_port, Q => err_1_port);
   err_reg_0_inst : DFFSR port map( D => n540, CLK => clk, R => n24, S => 
                           n108_port, Q => err_0_port);
   steep_reg : DFFSR port map( D => n539, CLK => clk, R => n24, S => n107_port,
                           Q => steep);
   Y_reg_0_inst : DFFSR port map( D => n518, CLK => clk, R => n24, S => 
                           n106_port, Q => N213);
   X_reg_0_inst : DFFSR port map( D => n510, CLK => clk, R => n24, S => 
                           n105_port, Q => N229);
   X_reg_7_inst : DFFSR port map( D => n499, CLK => clk, R => n24, S => 
                           n104_port, Q => N212);
   Y_reg_7_inst : DFFSR port map( D => n511, CLK => clk, R => n24, S => 
                           n103_port, Q => N220);
   Y_reg_6_inst : DFFSR port map( D => n512, CLK => clk, R => n24, S => 
                           n102_port, Q => N219);
   X_reg_6_inst : DFFSR port map( D => n500, CLK => clk, R => n24, S => 
                           n101_port, Q => N211);
   X_reg_5_inst : DFFSR port map( D => n501, CLK => clk, R => n25, S => 
                           n100_port, Q => N210);
   Y_reg_5_inst : DFFSR port map( D => n513, CLK => clk, R => n25, S => 
                           n99_port, Q => N218);
   Y_reg_1_inst : DFFSR port map( D => n517, CLK => clk, R => n25, S => 
                           n98_port, Q => N214);
   X_reg_1_inst : DFFSR port map( D => n509, CLK => clk, R => n25, S => 
                           n97_port, Q => N230);
   rast_indexi_reg_1_inst : DFFSR port map( D => n505, CLK => clk, R => n25, S 
                           => n96, Q => rast_index_1_port);
   Y_reg_2_inst : DFFSR port map( D => n516, CLK => clk, R => n25, S => 
                           n95_port, Q => N215);
   X_reg_2_inst : DFFSR port map( D => n508, CLK => clk, R => n25, S => n94, Q 
                           => N231);
   rast_indexi_reg_2_inst : DFFSR port map( D => n504, CLK => clk, R => n25, S 
                           => n93, Q => rast_index_2_port);
   Y_reg_3_inst : DFFSR port map( D => n515, CLK => clk, R => n25, S => n92, Q 
                           => N216);
   X_reg_3_inst : DFFSR port map( D => n507, CLK => clk, R => n25, S => n91, Q 
                           => N232);
   rast_indexi_reg_3_inst : DFFSR port map( D => n503, CLK => clk, R => n25, S 
                           => n90, Q => rast_index_3_port);
   Y_reg_4_inst : DFFSR port map( D => n514, CLK => clk, R => n26, S => n89, Q 
                           => N217);
   X_reg_4_inst : DFFSR port map( D => n502, CLK => clk, R => n26, S => n88, Q 
                           => N209);
   rast_addri_reg_4_inst : DFFSR port map( D => n498, CLK => clk, R => n26, S 
                           => n87, Q => rast_addr_0_port);
   rast_addri_reg_5_inst : DFFSR port map( D => n497, CLK => clk, R => n26, S 
                           => n86, Q => rast_addr_1_port);
   rast_addri_reg_6_inst : DFFSR port map( D => n496, CLK => clk, R => n25, S 
                           => n85, Q => rast_addr_2_port);
   rast_addri_reg_7_inst : DFFSR port map( D => n495, CLK => clk, R => n26, S 
                           => n84, Q => rast_addr_3_port);
   rast_addri_reg_8_inst : DFFSR port map( D => n494, CLK => clk, R => n26, S 
                           => n83, Q => rast_addr_4_port);
   rast_addri_reg_9_inst : DFFSR port map( D => n493, CLK => clk, R => n26, S 
                           => n82, Q => rast_addr_5_port);
   rast_addri_reg_10_inst : DFFSR port map( D => n492, CLK => clk, R => n26, S 
                           => n81, Q => rast_addr_6_port);
   rast_addri_reg_11_inst : DFFSR port map( D => n491, CLK => clk, R => n26, S 
                           => n80, Q => rast_addr_7_port);
   rast_addri_reg_12_inst : DFFSR port map( D => n490, CLK => clk, R => n26, S 
                           => n79, Q => rast_addr_8_port);
   rast_addri_reg_13_inst : DFFSR port map( D => n489, CLK => clk, R => n26, S 
                           => n78, Q => rast_addr_9_port);
   rast_addri_reg_14_inst : DFFSR port map( D => n488, CLK => clk, R => n26, S 
                           => n77, Q => rast_addr_10_port);
   rast_addri_reg_15_inst : DFFSR port map( D => n487, CLK => clk, R => n27, S 
                           => n76, Q => rast_addr_11_port);
   rast_indexi_reg_0_inst : DFFSR port map( D => n506, CLK => clk, R => n27, S 
                           => n75, Q => rast_index_0_port);
   i_reg_7_inst : DFFSR port map( D => n568, CLK => clk, R => n27, S => n74, Q 
                           => i_7_port);
   i_reg_1_inst : DFFSR port map( D => n574, CLK => clk, R => n27, S => n73, Q 
                           => i_1_port);
   i_reg_2_inst : DFFSR port map( D => n573, CLK => clk, R => n27, S => n72, Q 
                           => i_2_port);
   i_reg_3_inst : DFFSR port map( D => n572, CLK => clk, R => n27, S => n71, Q 
                           => i_3_port);
   i_reg_4_inst : DFFSR port map( D => n571, CLK => clk, R => n27, S => n70, Q 
                           => i_4_port);
   i_reg_5_inst : DFFSR port map( D => n570, CLK => clk, R => n27, S => n69, Q 
                           => i_5_port);
   i_reg_6_inst : DFFSR port map( D => n569, CLK => clk, R => n21, S => n68, Q 
                           => i_6_port);
   n68 <= '1';
   n69 <= '1';
   n70 <= '1';
   n71 <= '1';
   n72 <= '1';
   n73 <= '1';
   n74 <= '1';
   n75 <= '1';
   n76 <= '1';
   n77 <= '1';
   n78 <= '1';
   n79 <= '1';
   n80 <= '1';
   n81 <= '1';
   n82 <= '1';
   n83 <= '1';
   n84 <= '1';
   n85 <= '1';
   n86 <= '1';
   n87 <= '1';
   n88 <= '1';
   n89 <= '1';
   n90 <= '1';
   n91 <= '1';
   n92 <= '1';
   n93 <= '1';
   n94 <= '1';
   n95_port <= '1';
   n96 <= '1';
   n97_port <= '1';
   n98_port <= '1';
   n99_port <= '1';
   n100_port <= '1';
   n101_port <= '1';
   n102_port <= '1';
   n103_port <= '1';
   n104_port <= '1';
   n105_port <= '1';
   n106_port <= '1';
   n107_port <= '1';
   n108_port <= '1';
   n109_port <= '1';
   n110_port <= '1';
   n111_port <= '1';
   n112_port <= '1';
   n113 <= '1';
   n114 <= '1';
   n115 <= '1';
   n116 <= '1';
   n117 <= '1';
   n118 <= '1';
   n119 <= '1';
   n120 <= '1';
   n121_port <= '1';
   n122 <= '1';
   n123_port <= '1';
   n124_port <= '1';
   n125_port <= '1';
   n126_port <= '1';
   n127_port <= '1';
   n128_port <= '1';
   n129_port <= '1';
   n130_port <= '1';
   n131_port <= '1';
   n132_port <= '1';
   n133_port <= '1';
   n134_port <= '1';
   n135_port <= '1';
   n136_port <= '1';
   n137_port <= '1';
   n138_port <= '1';
   n139 <= '1';
   n140 <= '1';
   n141 <= '1';
   n142 <= '1';
   n143 <= '1';
   n144 <= '1';
   n145 <= '1';
   n146 <= '1';
   n147 <= '1';
   n148 <= '1';
   U102 : AND2X2 port map( A => n255, B => n256, Y => n249);
   U104 : OR2X2 port map( A => n312_port, B => n612, Y => n281_port);
   U105 : OR2X2 port map( A => n312_port, B => n611, Y => n317_port);
   U106 : AND2X2 port map( A => state_1_port, B => n616, Y => n477);
   U107 : AND2X2 port map( A => state_1_port, B => state_0_port, Y => n484);
   U188 : NOR2X1 port map( A => n229_port, B => n230_port, Y => rast_strb);
   U189 : NAND2X1 port map( A => n599, B => n621, Y => n230_port);
   U190 : NAND3X1 port map( A => n623, B => n618, C => n622, Y => n229_port);
   U191 : NAND3X1 port map( A => n598, B => n231_port, C => n232_port, Y => 
                           nextstate_3_port);
   U192 : NOR2X1 port map( A => n612, B => n233, Y => n232_port);
   U193 : NAND2X1 port map( A => n234, B => n235, Y => n233);
   U194 : OAI21X1 port map( A => count_2_port, B => n236, C => n599, Y => 
                           n231_port);
   U195 : NAND3X1 port map( A => n237, B => n598, C => n238, Y => 
                           nextstate_2_port);
   U196 : NOR2X1 port map( A => n239, B => n240, Y => n238);
   U197 : NAND2X1 port map( A => n241, B => n242, Y => n240);
   U198 : NAND2X1 port map( A => n243, B => n244, Y => n239);
   U199 : OAI21X1 port map( A => n246, B => n247, C => n248, Y => n245);
   U200 : NOR2X1 port map( A => n236, B => n623, Y => n246);
   U201 : AOI21X1 port map( A => N265, B => n601, C => n611, Y => n237);
   U202 : NAND3X1 port map( A => n249, B => n250, C => n251, Y => 
                           nextstate_1_port);
   U203 : NOR2X1 port map( A => n610, B => n252, Y => n251);
   U204 : OAI21X1 port map( A => N266, B => n234, C => n253, Y => n252);
   U205 : NAND3X1 port map( A => n599, B => n623, C => n617, Y => n253);
   U206 : NAND3X1 port map( A => n622, B => n618, C => count_0_port, Y => n236)
                           ;
   U207 : NOR2X1 port map( A => n603, B => n606, Y => n250);
   U208 : NAND3X1 port map( A => n257_port, B => n258_port, C => n259_port, Y 
                           => nextstate_0_port);
   U209 : NOR2X1 port map( A => n260_port, B => n261_port, Y => n259_port);
   U210 : NAND2X1 port map( A => n262_port, B => n243, Y => n261_port);
   U211 : NAND2X1 port map( A => n248, B => n244, Y => n260_port);
   U212 : AOI21X1 port map( A => init_rast, B => n608, C => n605, Y => 
                           n258_port);
   U213 : AOI22X1 port map( A => N266, B => n609, C => n607, D => n613, Y => 
                           n257_port);
   U214 : OAI21X1 port map( A => n576, B => n641, C => n263_port, Y => n487);
   U215 : AOI22X1 port map( A => N220, B => n9, C => N212, D => n1, Y => 
                           n263_port);
   U216 : OAI21X1 port map( A => n576, B => n640, C => n266_port, Y => n488);
   U217 : AOI22X1 port map( A => N219, B => n9, C => N211, D => n1, Y => 
                           n266_port);
   U218 : OAI21X1 port map( A => n576, B => n639, C => n267, Y => n489);
   U219 : AOI22X1 port map( A => N218, B => n9, C => N210, D => n1, Y => n267);
   U220 : OAI21X1 port map( A => n576, B => n638, C => n268, Y => n490);
   U221 : AOI22X1 port map( A => N217, B => n9, C => N209, D => n1, Y => n268);
   U222 : OAI21X1 port map( A => n576, B => n637, C => n269_port, Y => n491);
   U223 : AOI22X1 port map( A => N216, B => n9, C => N232, D => n1, Y => 
                           n269_port);
   U224 : OAI21X1 port map( A => n576, B => n636, C => n270_port, Y => n492);
   U225 : AOI22X1 port map( A => N215, B => n9, C => N231, D => n1, Y => 
                           n270_port);
   U226 : OAI21X1 port map( A => n576, B => n635, C => n271_port, Y => n493);
   U227 : AOI22X1 port map( A => N214, B => n9, C => N230, D => n1, Y => 
                           n271_port);
   U228 : OAI21X1 port map( A => n576, B => n634, C => n272_port, Y => n494);
   U229 : AOI22X1 port map( A => N213, B => n9, C => N229, D => n1, Y => 
                           n272_port);
   U230 : OAI21X1 port map( A => n576, B => n633, C => n273_port, Y => n495);
   U231 : AOI22X1 port map( A => N212, B => n9, C => N220, D => n1, Y => 
                           n273_port);
   U232 : OAI21X1 port map( A => n576, B => n632, C => n274_port, Y => n496);
   U233 : AOI22X1 port map( A => N211, B => n9, C => N219, D => n1, Y => 
                           n274_port);
   U234 : OAI21X1 port map( A => n576, B => n631, C => n275_port, Y => n497);
   U235 : AOI22X1 port map( A => N210, B => n9, C => N218, D => n1, Y => 
                           n275_port);
   U236 : OAI21X1 port map( A => n576, B => n630, C => n276_port, Y => n498);
   U237 : AOI22X1 port map( A => N209, B => n9, C => N217, D => n1, Y => 
                           n276_port);
   U238 : NAND3X1 port map( A => n277_port, B => n278_port, C => n279_port, Y 
                           => n499);
   U239 : AOI22X1 port map( A => N333, B => n280_port, C => N212, D => 
                           n281_port, Y => n279_port);
   U240 : NAND2X1 port map( A => N325, B => n282_port, Y => n278_port);
   U241 : AOI22X1 port map( A => N220, B => n283_port, C => X0(7), D => n606, Y
                           => n277_port);
   U242 : NAND3X1 port map( A => n284_port, B => n285_port, C => n286_port, Y 
                           => n500);
   U243 : AOI22X1 port map( A => N332, B => n280_port, C => N211, D => 
                           n281_port, Y => n286_port);
   U244 : NAND2X1 port map( A => N324, B => n282_port, Y => n285_port);
   U245 : AOI22X1 port map( A => N219, B => n283_port, C => X0(6), D => n606, Y
                           => n284_port);
   U246 : NAND3X1 port map( A => n287_port, B => n288_port, C => n289_port, Y 
                           => n501);
   U247 : AOI22X1 port map( A => N331, B => n280_port, C => N210, D => 
                           n281_port, Y => n289_port);
   U248 : NAND2X1 port map( A => N323, B => n282_port, Y => n288_port);
   U249 : AOI22X1 port map( A => N218, B => n283_port, C => X0(5), D => n606, Y
                           => n287_port);
   U250 : NAND3X1 port map( A => n290_port, B => n291_port, C => n292_port, Y 
                           => n502);
   U251 : AOI22X1 port map( A => N330, B => n280_port, C => N209, D => 
                           n281_port, Y => n292_port);
   U252 : NAND2X1 port map( A => N322, B => n282_port, Y => n291_port);
   U253 : AOI22X1 port map( A => N217, B => n283_port, C => X0(4), D => n606, Y
                           => n290_port);
   U254 : OAI21X1 port map( A => n576, B => n629, C => n293_port, Y => n503);
   U255 : AOI22X1 port map( A => N232, B => n9, C => N216, D => n1, Y => 
                           n293_port);
   U256 : OAI21X1 port map( A => n576, B => n628, C => n294_port, Y => n504);
   U257 : AOI22X1 port map( A => N231, B => n9, C => N215, D => n1, Y => 
                           n294_port);
   U258 : OAI21X1 port map( A => n576, B => n627, C => n295_port, Y => n505);
   U259 : AOI22X1 port map( A => N230, B => n9, C => N214, D => n1, Y => 
                           n295_port);
   U260 : OAI21X1 port map( A => n576, B => n642, C => n296_port, Y => n506);
   U261 : AOI22X1 port map( A => N229, B => n9, C => N213, D => n1, Y => 
                           n296_port);
   U263 : NAND3X1 port map( A => n298, B => n235, C => n577, Y => n297);
   U264 : NAND3X1 port map( A => n299, B => n300, C => n301, Y => n507);
   U265 : AOI22X1 port map( A => N329, B => n280_port, C => N232, D => 
                           n281_port, Y => n301);
   U266 : NAND2X1 port map( A => N321, B => n282_port, Y => n300);
   U267 : AOI22X1 port map( A => N216, B => n283_port, C => X0(3), D => n606, Y
                           => n299);
   U268 : NAND3X1 port map( A => n302, B => n303, C => n304, Y => n508);
   U269 : AOI22X1 port map( A => N328, B => n280_port, C => N231, D => 
                           n281_port, Y => n304);
   U270 : NAND2X1 port map( A => N320, B => n282_port, Y => n303);
   U271 : AOI22X1 port map( A => N215, B => n283_port, C => X0(2), D => n606, Y
                           => n302);
   U272 : NAND3X1 port map( A => n305, B => n306_port, C => n307_port, Y => 
                           n509);
   U273 : AOI22X1 port map( A => N327, B => n280_port, C => N230, D => 
                           n281_port, Y => n307_port);
   U274 : NAND2X1 port map( A => N319, B => n282_port, Y => n306_port);
   U275 : AOI22X1 port map( A => N214, B => n283_port, C => X0(1), D => n606, Y
                           => n305);
   U276 : NAND3X1 port map( A => n308_port, B => n309_port, C => n310_port, Y 
                           => n510);
   U277 : AOI22X1 port map( A => N326, B => n280_port, C => N229, D => 
                           n281_port, Y => n310_port);
   U278 : NOR2X1 port map( A => n624, B => n311_port, Y => n280_port);
   U279 : NAND2X1 port map( A => N318, B => n282_port, Y => n309_port);
   U280 : NOR2X1 port map( A => n311_port, B => iX, Y => n282_port);
   U281 : AOI22X1 port map( A => N213, B => n283_port, C => X0(0), D => n606, Y
                           => n308_port);
   U282 : NOR2X1 port map( A => n281_port, B => n243, Y => n283_port);
   U283 : NAND3X1 port map( A => n313_port, B => n314_port, C => n315_port, Y 
                           => n511);
   U284 : AOI22X1 port map( A => N296, B => n316_port, C => N220, D => 
                           n317_port, Y => n315_port);
   U285 : NAND2X1 port map( A => N288, B => n318_port, Y => n314_port);
   U286 : AOI22X1 port map( A => n319_port, B => N212, C => Y0(7), D => n606, Y
                           => n313_port);
   U287 : NAND3X1 port map( A => n320_port, B => n321_port, C => n322_port, Y 
                           => n512);
   U288 : AOI22X1 port map( A => N295, B => n316_port, C => N219, D => 
                           n317_port, Y => n322_port);
   U289 : NAND2X1 port map( A => N287, B => n318_port, Y => n321_port);
   U290 : AOI22X1 port map( A => n319_port, B => N211, C => Y0(6), D => n606, Y
                           => n320_port);
   U291 : NAND3X1 port map( A => n323_port, B => n324_port, C => n325_port, Y 
                           => n513);
   U292 : AOI22X1 port map( A => N294, B => n316_port, C => N218, D => 
                           n317_port, Y => n325_port);
   U293 : NAND2X1 port map( A => N286, B => n318_port, Y => n324_port);
   U294 : AOI22X1 port map( A => n319_port, B => N210, C => Y0(5), D => n606, Y
                           => n323_port);
   U295 : NAND3X1 port map( A => n326_port, B => n327_port, C => n328_port, Y 
                           => n514);
   U296 : AOI22X1 port map( A => N293, B => n316_port, C => N217, D => 
                           n317_port, Y => n328_port);
   U297 : NAND2X1 port map( A => N285, B => n318_port, Y => n327_port);
   U298 : AOI22X1 port map( A => n319_port, B => N209, C => Y0(4), D => n606, Y
                           => n326_port);
   U299 : NAND3X1 port map( A => n329_port, B => n330_port, C => n331_port, Y 
                           => n515);
   U300 : AOI22X1 port map( A => N292, B => n316_port, C => N216, D => 
                           n317_port, Y => n331_port);
   U301 : NAND2X1 port map( A => N284, B => n318_port, Y => n330_port);
   U302 : AOI22X1 port map( A => n319_port, B => N232, C => Y0(3), D => n606, Y
                           => n329_port);
   U303 : NAND3X1 port map( A => n332_port, B => n333_port, C => n334, Y => 
                           n516);
   U304 : AOI22X1 port map( A => N291, B => n316_port, C => N215, D => 
                           n317_port, Y => n334);
   U305 : NAND2X1 port map( A => N283, B => n318_port, Y => n333_port);
   U306 : AOI22X1 port map( A => n319_port, B => N231, C => Y0(2), D => n606, Y
                           => n332_port);
   U307 : NAND3X1 port map( A => n335, B => n336, C => n337, Y => n517);
   U308 : AOI22X1 port map( A => N290, B => n316_port, C => N214, D => 
                           n317_port, Y => n337);
   U309 : NAND2X1 port map( A => N282, B => n318_port, Y => n336);
   U310 : AOI22X1 port map( A => n319_port, B => N230, C => Y0(1), D => n606, Y
                           => n335);
   U311 : NAND3X1 port map( A => n338, B => n339, C => n340, Y => n518);
   U312 : AOI22X1 port map( A => N289, B => n316_port, C => N213, D => 
                           n317_port, Y => n340);
   U313 : NOR2X1 port map( A => n625, B => n341, Y => n316_port);
   U314 : NAND2X1 port map( A => N281, B => n318_port, Y => n339);
   U315 : NOR2X1 port map( A => n341, B => iY, Y => n318_port);
   U316 : AOI22X1 port map( A => n319_port, B => N229, C => Y0(0), D => n606, Y
                           => n338);
   U317 : NOR2X1 port map( A => n317_port, B => n243, Y => n319_port);
   U318 : NAND3X1 port map( A => n342, B => n298, C => n343, Y => n312_port);
   U319 : NOR2X1 port map( A => n607, B => n605, Y => n343);
   U320 : OAI21X1 port map( A => n594, B => n624, C => n344, Y => n519);
   U321 : OAI21X1 port map( A => n345, B => n346, C => n594, Y => n344);
   U323 : OAI21X1 port map( A => n594, B => n625, C => n347, Y => n520);
   U324 : OAI21X1 port map( A => n348, B => n349, C => n594, Y => n347);
   U326 : NAND3X1 port map( A => n254, B => n242, C => n342, Y => n350);
   U327 : AOI22X1 port map( A => N264, B => n601, C => i_7_port, D => n352, Y 
                           => n351);
   U328 : AOI22X1 port map( A => N263, B => n601, C => i_6_port, D => n352, Y 
                           => n353);
   U329 : AOI22X1 port map( A => N262, B => n601, C => i_5_port, D => n352, Y 
                           => n354);
   U330 : AOI22X1 port map( A => N261, B => n601, C => i_4_port, D => n352, Y 
                           => n355);
   U331 : AOI22X1 port map( A => N260, B => n601, C => i_3_port, D => n352, Y 
                           => n356);
   U332 : AOI22X1 port map( A => N259, B => n601, C => i_2_port, D => n352, Y 
                           => n357);
   U333 : AOI22X1 port map( A => N258, B => n601, C => i_1_port, D => n352, Y 
                           => n358);
   U334 : NAND2X1 port map( A => n359, B => n360, Y => n521);
   U336 : AOI22X1 port map( A => dy_8_port, B => n8, C => dx_8_port, D => n7, Y
                           => n359);
   U337 : NAND3X1 port map( A => n364, B => n365, C => n366, Y => n522);
   U338 : AOI21X1 port map( A => n10, B => n7, C => n593, Y => n366);
   U339 : AOI22X1 port map( A => n8, B => dy_7_port, C => n607, D => n11, Y => 
                           n367);
   U340 : NAND2X1 port map( A => N104, B => n345, Y => n365);
   U342 : NAND3X1 port map( A => n369, B => n370, C => n371, Y => n523);
   U343 : AOI21X1 port map( A => n11, B => n7, C => n592, Y => n371);
   U344 : AOI22X1 port map( A => n8, B => dy_6_port, C => n607, D => n12, Y => 
                           n372);
   U345 : NAND2X1 port map( A => N103, B => n345, Y => n370);
   U347 : NAND3X1 port map( A => n373, B => n374, C => n375, Y => n524);
   U348 : AOI21X1 port map( A => n12, B => n7, C => n591, Y => n375);
   U349 : AOI22X1 port map( A => n8, B => dy_5_port, C => n607, D => n15, Y => 
                           n376);
   U350 : NAND2X1 port map( A => N102, B => n345, Y => n374);
   U352 : NAND3X1 port map( A => n377, B => n378, C => n379, Y => n525);
   U353 : AOI21X1 port map( A => n15, B => n7, C => n590, Y => n379);
   U354 : AOI22X1 port map( A => n8, B => dy_4_port, C => n607, D => n18, Y => 
                           n380);
   U355 : NAND2X1 port map( A => N101, B => n345, Y => n378);
   U357 : NAND3X1 port map( A => n381, B => n382, C => n383, Y => n526);
   U358 : AOI21X1 port map( A => n18, B => n7, C => n589, Y => n383);
   U359 : AOI22X1 port map( A => n8, B => dy_3_port, C => n607, D => n19, Y => 
                           n384);
   U360 : NAND2X1 port map( A => N100, B => n345, Y => n382);
   U362 : NAND3X1 port map( A => n385, B => n386, C => n387, Y => n527);
   U363 : AOI21X1 port map( A => n19, B => n7, C => n588, Y => n387);
   U364 : AOI22X1 port map( A => n8, B => dy_2_port, C => n607, D => N190, Y =>
                           n388);
   U365 : NAND2X1 port map( A => N99, B => n345, Y => n386);
   U367 : NAND3X1 port map( A => n389, B => n390, C => n391, Y => n528);
   U368 : AOI21X1 port map( A => N190, B => n7, C => n587, Y => n391);
   U369 : AOI22X1 port map( A => n8, B => dy_1_port, C => n607, D => dx_0_port,
                           Y => n392);
   U370 : NAND2X1 port map( A => N98, B => n345, Y => n390);
   U372 : NAND3X1 port map( A => n393, B => n394, C => n395, Y => n529);
   U373 : AOI22X1 port map( A => dy_0_port, B => n8, C => dx_0_port, D => n7, Y
                           => n395);
   U375 : NAND2X1 port map( A => N97, B => n345, Y => n394);
   U376 : NOR2X1 port map( A => n566, B => n262_port, Y => n345);
   U378 : NOR2X1 port map( A => n262_port, B => N95, Y => n368);
   U380 : NAND2X1 port map( A => n396, B => n397, Y => n530);
   U382 : AOI22X1 port map( A => dx_8_port, B => n8, C => dy_8_port, D => n363,
                           Y => n396);
   U383 : NAND3X1 port map( A => n400, B => n401, C => n402, Y => n531);
   U384 : AOI21X1 port map( A => dy_7_port, B => n363, C => n586, Y => n402);
   U385 : AOI22X1 port map( A => n10, B => n8, C => n607, D => dy_6_port, Y => 
                           n403);
   U386 : NAND2X1 port map( A => N130, B => n348, Y => n401);
   U388 : NAND3X1 port map( A => n405, B => n406, C => n407, Y => n532);
   U389 : AOI21X1 port map( A => dy_6_port, B => n363, C => n585, Y => n407);
   U390 : AOI22X1 port map( A => n8, B => n11, C => n607, D => dy_5_port, Y => 
                           n408);
   U391 : NAND2X1 port map( A => N129, B => n348, Y => n406);
   U393 : NAND3X1 port map( A => n409, B => n410, C => n411, Y => n533);
   U394 : AOI21X1 port map( A => dy_5_port, B => n363, C => n584, Y => n411);
   U395 : AOI22X1 port map( A => n8, B => n12, C => n607, D => dy_4_port, Y => 
                           n412);
   U396 : NAND2X1 port map( A => N128, B => n348, Y => n410);
   U398 : NAND3X1 port map( A => n413, B => n414, C => n415, Y => n534);
   U399 : AOI21X1 port map( A => dy_4_port, B => n363, C => n583, Y => n415);
   U400 : AOI22X1 port map( A => n8, B => n15, C => n607, D => dy_3_port, Y => 
                           n416);
   U401 : NAND2X1 port map( A => N127, B => n348, Y => n414);
   U403 : NAND3X1 port map( A => n417, B => n418, C => n419, Y => n535);
   U404 : AOI21X1 port map( A => dy_3_port, B => n363, C => n582, Y => n419);
   U405 : AOI22X1 port map( A => n8, B => n18, C => n607, D => dy_2_port, Y => 
                           n420);
   U406 : NAND2X1 port map( A => N126, B => n348, Y => n418);
   U408 : NAND3X1 port map( A => n421, B => n422, C => n423, Y => n536);
   U409 : AOI21X1 port map( A => dy_2_port, B => n363, C => n581, Y => n423);
   U410 : AOI22X1 port map( A => n8, B => n19, C => n607, D => dy_1_port, Y => 
                           n424);
   U411 : NAND2X1 port map( A => N125, B => n348, Y => n422);
   U413 : NAND3X1 port map( A => n425, B => n426, C => n427, Y => n537);
   U414 : AOI21X1 port map( A => dy_1_port, B => n363, C => n580, Y => n427);
   U415 : AOI22X1 port map( A => n8, B => N190, C => n607, D => dy_0_port, Y =>
                           n428);
   U416 : NAND2X1 port map( A => N124, B => n348, Y => n426);
   U418 : NAND3X1 port map( A => n429, B => n430, C => n431, Y => n538);
   U419 : AOI22X1 port map( A => dx_0_port, B => n8, C => dy_0_port, D => n363,
                           Y => n431);
   U422 : NAND3X1 port map( A => n254, B => n298, C => n342, Y => n432);
   U423 : NOR3X1 port map( A => n603, B => n609, C => n433, Y => n342);
   U424 : OAI21X1 port map( A => n243, B => steep, C => n595, Y => n433);
   U425 : NAND2X1 port map( A => N123, B => n348, Y => n430);
   U426 : NOR2X1 port map( A => n565, B => n262_port, Y => n348);
   U428 : NOR2X1 port map( A => n262_port, B => N121, Y => n404);
   U430 : OAI21X1 port map( A => n242, B => n613, C => n434, Y => n539);
   U431 : OAI21X1 port map( A => n602, B => n435, C => steep, Y => n434);
   U432 : NAND2X1 port map( A => n437, B => n438, Y => n540);
   U433 : AOI22X1 port map( A => N199, B => n603, C => N306, D => n611, Y => 
                           n438);
   U434 : AOI22X1 port map( A => N269, B => n612, C => err_0_port, D => n578, Y
                           => n437);
   U435 : NAND2X1 port map( A => n439, B => n440, Y => n541);
   U436 : AOI22X1 port map( A => N200, B => n603, C => N307, D => n611, Y => 
                           n440);
   U437 : AOI22X1 port map( A => N270, B => n612, C => err_1_port, D => n578, Y
                           => n439);
   U438 : NAND2X1 port map( A => n441, B => n442, Y => n542);
   U439 : AOI22X1 port map( A => N201, B => n603, C => N308, D => n611, Y => 
                           n442);
   U440 : AOI22X1 port map( A => N271, B => n612, C => err_2_port, D => n578, Y
                           => n441);
   U441 : NAND2X1 port map( A => n443, B => n444, Y => n543);
   U442 : AOI22X1 port map( A => N202, B => n603, C => N309, D => n611, Y => 
                           n444);
   U443 : AOI22X1 port map( A => N272, B => n612, C => err_3_port, D => n578, Y
                           => n443);
   U444 : NAND2X1 port map( A => n445, B => n446, Y => n544);
   U445 : AOI22X1 port map( A => N203, B => n603, C => N310, D => n611, Y => 
                           n446);
   U446 : AOI22X1 port map( A => N273, B => n612, C => err_4_port, D => n578, Y
                           => n445);
   U447 : NAND2X1 port map( A => n447, B => n448, Y => n545);
   U448 : AOI22X1 port map( A => N204, B => n603, C => N311, D => n611, Y => 
                           n448);
   U449 : AOI22X1 port map( A => N274, B => n612, C => err_5_port, D => n578, Y
                           => n447);
   U450 : NAND2X1 port map( A => n449, B => n450, Y => n546);
   U451 : AOI22X1 port map( A => N205, B => n603, C => N312, D => n611, Y => 
                           n450);
   U452 : AOI22X1 port map( A => N275, B => n612, C => err_6_port, D => n578, Y
                           => n449);
   U453 : NAND2X1 port map( A => n451, B => n452, Y => n547);
   U454 : AOI22X1 port map( A => N206, B => n603, C => N313, D => n611, Y => 
                           n452);
   U455 : AOI22X1 port map( A => N276, B => n612, C => err_7_port, D => n578, Y
                           => n451);
   U456 : OAI21X1 port map( A => n453, B => n626, C => n454, Y => n548);
   U457 : AOI22X1 port map( A => N315, B => n611, C => N278, D => n612, Y => 
                           n454);
   U458 : OAI21X1 port map( A => n453, B => n615, C => n455, Y => n549);
   U459 : AOI22X1 port map( A => N316, B => n611, C => N279, D => n612, Y => 
                           n455);
   U460 : OAI22X1 port map( A => n600, B => n618, C => n456, D => n457, Y => 
                           n550);
   U461 : XNOR2X1 port map( A => count_3_port, B => n458, Y => n457);
   U462 : NOR2X1 port map( A => n623, B => n620, Y => n458);
   U463 : OAI21X1 port map( A => n459, B => n623, C => n460, Y => n551);
   U464 : NAND3X1 port map( A => n575, B => n623, C => n461, Y => n460);
   U465 : AOI21X1 port map( A => n620, B => n575, C => n462, Y => n459);
   U466 : NOR2X1 port map( A => n622, B => n621, Y => n461);
   U467 : OAI21X1 port map( A => n463, B => n622, C => n464, Y => n552);
   U468 : NAND3X1 port map( A => n575, B => n622, C => count_0_port, Y => n464)
                           ;
   U469 : AOI21X1 port map( A => n575, B => n621, C => n462, Y => n463);
   U470 : OAI22X1 port map( A => n600, B => n621, C => count_0_port, D => n456,
                           Y => n553);
   U471 : NAND3X1 port map( A => n436, B => n465, C => n466, Y => n462);
   U472 : NOR2X1 port map( A => n608, B => n467, Y => n466);
   U473 : NAND2X1 port map( A => n256, B => n242, Y => n467);
   U474 : OAI21X1 port map( A => n453, B => n614, C => n468, Y => n554);
   U475 : AOI22X1 port map( A => N317, B => n611, C => N280, D => n612, Y => 
                           n468);
   U476 : NAND3X1 port map( A => n469, B => n470, C => n471, Y => n555);
   U477 : AOI21X1 port map( A => err_8_port, B => n578, C => n608, Y => n471);
   U478 : NAND2X1 port map( A => n472, B => n473, Y => n298);
   U479 : NOR2X1 port map( A => n474, B => n475, Y => n453);
   U480 : NAND3X1 port map( A => n255, B => n262_port, C => n595, Y => n475);
   U481 : NAND3X1 port map( A => n248, B => n235, C => n596, Y => n435);
   U482 : NAND3X1 port map( A => n243, B => n234, C => n242, Y => n474);
   U483 : NAND2X1 port map( A => N277, B => n612, Y => n470);
   U484 : AOI22X1 port map( A => N207, B => n603, C => N314, D => n611, Y => 
                           n469);
   U485 : AOI22X1 port map( A => N257, B => n601, C => i_0_port, D => n352, Y 
                           => n476);
   U486 : NAND2X1 port map( A => n577, B => n248, Y => n352);
   U487 : NAND2X1 port map( A => n477, B => n478, Y => n248);
   U488 : NAND3X1 port map( A => n436, B => n242, C => n596, Y => n479);
   U489 : NAND3X1 port map( A => n256, B => n456, C => n465, Y => n480);
   U490 : NAND2X1 port map( A => state_1_port, B => n481, Y => n465);
   U491 : NOR2X1 port map( A => rast_done_port, B => n599, Y => n456);
   U492 : NAND2X1 port map( A => n481, B => n482, Y => n244);
   U493 : NAND2X1 port map( A => n483, B => n484, Y => n256);
   U494 : NAND2X1 port map( A => n472, B => n484, Y => n242);
   U495 : NOR2X1 port map( A => n485, B => n486, Y => n436);
   U496 : NAND3X1 port map( A => n255, B => n262_port, C => n254, Y => n486);
   U497 : NOR2X1 port map( A => n611, B => n612, Y => n254);
   U498 : NAND2X1 port map( A => n483, B => n482, Y => n341);
   U499 : NAND2X1 port map( A => n477, B => n483, Y => n311_port);
   U500 : NAND2X1 port map( A => n472, B => n482, Y => n262_port);
   U501 : NAND2X1 port map( A => n472, B => n477, Y => n255);
   U502 : NOR2X1 port map( A => state_2_port, B => state_3_port, Y => n472);
   U503 : NAND3X1 port map( A => n243, B => n234, C => n241, Y => n485);
   U504 : NAND2X1 port map( A => n478, B => n482, Y => n241);
   U505 : NOR2X1 port map( A => n616, B => state_1_port, Y => n482);
   U506 : NAND2X1 port map( A => n473, B => n483, Y => n234);
   U507 : NOR2X1 port map( A => n619, B => state_2_port, Y => n483);
   U508 : NAND2X1 port map( A => n473, B => n478, Y => n243);
   U509 : NAND2X1 port map( A => n478, B => n484, Y => n235);
   U510 : NOR2X1 port map( A => n604, B => state_3_port, Y => n478);
   U511 : NAND2X1 port map( A => n473, B => n481, Y => n247);
   U512 : NOR2X1 port map( A => n619, B => n604, Y => n481);
   U513 : NOR2X1 port map( A => state_0_port, B => state_1_port, Y => n473);
   add_262 : Rasterizer_DW01_inc_0 port map( A(7) => N212, A(6) => N211, A(5) 
                           => N210, A(4) => N209, A(3) => N232, A(2) => N231, 
                           A(1) => N230, A(0) => N229, SUM(7) => N325, SUM(6) 
                           => N324, SUM(5) => N323, SUM(4) => N322, SUM(3) => 
                           N321, SUM(2) => N320, SUM(1) => N319, SUM(0) => N318
                           );
   add_259 : Rasterizer_DW01_add_0 port map( A(11) => err_11_port, A(10) => 
                           err_10_port, A(9) => err_9_port, A(8) => err_8_port,
                           A(7) => err_7_port, A(6) => err_6_port, A(5) => 
                           err_5_port, A(4) => err_4_port, A(3) => err_3_port, 
                           A(2) => err_2_port, A(1) => err_1_port, A(0) => 
                           err_0_port, B(11) => n3, B(10) => n3, B(9) => n3, 
                           B(8) => dy_8_port, B(7) => dy_7_port, B(6) => 
                           dy_6_port, B(5) => dy_5_port, B(4) => dy_4_port, 
                           B(3) => dy_3_port, B(2) => dy_2_port, B(1) => 
                           dy_1_port, B(0) => dy_0_port, CI => n3, SUM(11) => 
                           N317, SUM(10) => N316, SUM(9) => N315, SUM(8) => 
                           N314, SUM(7) => N313, SUM(6) => N312, SUM(5) => N311
                           , SUM(4) => N310, SUM(3) => N309, SUM(2) => N308, 
                           SUM(1) => N307, SUM(0) => N306, CO => n_1224);
   add_249 : Rasterizer_DW01_inc_1 port map( A(7) => N220, A(6) => N219, A(5) 
                           => N218, A(4) => N217, A(3) => N216, A(2) => N215, 
                           A(1) => N214, A(0) => N213, SUM(7) => N288, SUM(6) 
                           => N287, SUM(5) => N286, SUM(4) => N285, SUM(3) => 
                           N284, SUM(2) => N283, SUM(1) => N282, SUM(0) => N281
                           );
   sub_246 : Rasterizer_DW01_sub_2 port map( A(11) => err_11_port, A(10) => 
                           err_10_port, A(9) => err_9_port, A(8) => err_8_port,
                           A(7) => err_7_port, A(6) => err_6_port, A(5) => 
                           err_5_port, A(4) => err_4_port, A(3) => err_3_port, 
                           A(2) => err_2_port, A(1) => err_1_port, A(0) => 
                           err_0_port, B(11) => n4, B(10) => n4, B(9) => n4, 
                           B(8) => dx_8_port, B(7) => n10, B(6) => n11, B(5) =>
                           n12, B(4) => n15, B(3) => n18, B(2) => n19, B(1) => 
                           N190, B(0) => dx_0_port, CI => n4, DIFF(11) => N280,
                           DIFF(10) => N279, DIFF(9) => N278, DIFF(8) => N277, 
                           DIFF(7) => N276, DIFF(6) => N275, DIFF(5) => N274, 
                           DIFF(4) => N273, DIFF(3) => N272, DIFF(2) => N271, 
                           DIFF(1) => N270, DIFF(0) => N269, CO => n_1225);
   add_222 : Rasterizer_DW01_inc_2 port map( A(7) => i_7_port, A(6) => i_6_port
                           , A(5) => i_5_port, A(4) => i_4_port, A(3) => 
                           i_3_port, A(2) => i_2_port, A(1) => i_1_port, A(0) 
                           => i_0_port, SUM(7) => N264, SUM(6) => N263, SUM(5) 
                           => N262, SUM(4) => N261, SUM(3) => N260, SUM(2) => 
                           N259, SUM(1) => N258, SUM(0) => N257);
   sub_126 : Rasterizer_DW01_sub_3 port map( A(7) => Y1(7), A(6) => Y1(6), A(5)
                           => Y1(5), A(4) => Y1(4), A(3) => Y1(3), A(2) => 
                           Y1(2), A(1) => Y1(1), A(0) => Y1(0), B(7) => Y0(7), 
                           B(6) => Y0(6), B(5) => Y0(5), B(4) => Y0(4), B(3) =>
                           Y0(3), B(2) => Y0(2), B(1) => Y0(1), B(0) => Y0(0), 
                           CI => n13, DIFF(7) => N138, DIFF(6) => N137, DIFF(5)
                           => N136, DIFF(4) => N135, DIFF(3) => N134, DIFF(2) 
                           => N133, DIFF(1) => N132, DIFF(0) => N131, CO => 
                           n_1226);
   sub_123 : Rasterizer_DW01_sub_4 port map( A(7) => Y0(7), A(6) => Y0(6), A(5)
                           => Y0(5), A(4) => Y0(4), A(3) => Y0(3), A(2) => 
                           Y0(2), A(1) => Y0(1), A(0) => Y0(0), B(7) => Y1(7), 
                           B(6) => Y1(6), B(5) => Y1(5), B(4) => Y1(4), B(3) =>
                           Y1(3), B(2) => Y1(2), B(1) => Y1(1), B(0) => Y1(0), 
                           CI => n14, DIFF(7) => N130, DIFF(6) => N129, DIFF(5)
                           => N128, DIFF(4) => N127, DIFF(3) => N126, DIFF(2) 
                           => N125, DIFF(1) => N124, DIFF(0) => N123, CO => 
                           n_1227);
   sub_116 : Rasterizer_DW01_sub_5 port map( A(7) => X1(7), A(6) => X1(6), A(5)
                           => X1(5), A(4) => X1(4), A(3) => X1(3), A(2) => 
                           X1(2), A(1) => X1(1), A(0) => X1(0), B(7) => X0(7), 
                           B(6) => X0(6), B(5) => X0(5), B(4) => X0(4), B(3) =>
                           X0(3), B(2) => X0(2), B(1) => X0(1), B(0) => X0(0), 
                           CI => n16, DIFF(7) => N112, DIFF(6) => N111, DIFF(5)
                           => N110, DIFF(4) => N109, DIFF(3) => N108, DIFF(2) 
                           => N107, DIFF(1) => N106, DIFF(0) => N105, CO => 
                           n_1228);
   sub_111 : Rasterizer_DW01_sub_6 port map( A(7) => X0(7), A(6) => X0(6), A(5)
                           => X0(5), A(4) => X0(4), A(3) => X0(3), A(2) => 
                           X0(2), A(1) => X0(1), A(0) => X0(0), B(7) => X1(7), 
                           B(6) => X1(6), B(5) => X1(5), B(4) => X1(4), B(3) =>
                           X1(3), B(2) => X1(2), B(1) => X1(1), B(0) => X1(0), 
                           CI => n17, DIFF(7) => N104, DIFF(6) => N103, DIFF(5)
                           => N102, DIFF(4) => N101, DIFF(3) => N100, DIFF(2) 
                           => N99, DIFF(1) => N98, DIFF(0) => N97, CO => n_1229
                           );
   add_0_root_sub_0_root_sub_184 : Rasterizer_DW01_add_3 port map( A(8) => 
                           dy_8_port, A(7) => dy_7_port, A(6) => dy_6_port, 
                           A(5) => dy_5_port, A(4) => dy_4_port, A(3) => 
                           dy_3_port, A(2) => dy_2_port, A(1) => dy_1_port, 
                           A(0) => dy_0_port, B(8) => N198, B(7) => N197, B(6) 
                           => N196, B(5) => N195, B(4) => N194, B(3) => N193, 
                           B(2) => N192, B(1) => N191, B(0) => N190, CI => n643
                           , SUM(8) => N207, SUM(7) => N206, SUM(6) => N205, 
                           SUM(5) => N204, SUM(4) => N203, SUM(3) => N202, 
                           SUM(2) => N201, SUM(1) => N200, SUM(0) => N199, CO 
                           => n_1230);
   U13 : AND2X2 port map( A => steep, B => n576, Y => n1);
   U14 : INVX2 port map( A => n297, Y => n576);
   U17 : INVX2 port map( A => n2, Y => n8);
   U18 : INVX2 port map( A => n453, Y => n578);
   U19 : OR2X2 port map( A => n432, B => n243, Y => n2);
   U20 : INVX2 port map( A => n311_port, Y => n611);
   U21 : INVX2 port map( A => n341, Y => n612);
   U22 : INVX2 port map( A => n6, Y => n7);
   U23 : INVX2 port map( A => n363, Y => n6);
   U24 : INVX2 port map( A => n242, Y => n607);
   U27 : INVX2 port map( A => n241, Y => n603);
   U30 : INVX2 port map( A => n262_port, Y => n606);
   U103 : INVX2 port map( A => n235, Y => n601);
   U108 : INVX2 port map( A => n5, Y => n9);
   U109 : BUFX2 port map( A => dx_2_port, Y => n19);
   U110 : BUFX2 port map( A => dx_3_port, Y => n18);
   U111 : INVX2 port map( A => N190, Y => n20);
   U112 : OR2X2 port map( A => n297, B => steep, Y => n5);
   U113 : BUFX2 port map( A => dx_5_port, Y => n12);
   U114 : BUFX2 port map( A => dx_4_port, Y => n15);
   U115 : BUFX2 port map( A => dx_6_port, Y => n11);
   U116 : BUFX2 port map( A => dx_7_port, Y => n10);
   U117 : BUFX2 port map( A => RST_N, Y => n26);
   U118 : BUFX2 port map( A => RST_N, Y => n25);
   U119 : BUFX2 port map( A => RST_N, Y => n23);
   U120 : BUFX2 port map( A => RST_N, Y => n22);
   U121 : BUFX2 port map( A => RST_N, Y => n21);
   U122 : BUFX2 port map( A => RST_N, Y => n24);
   U123 : BUFX2 port map( A => RST_N, Y => n27);
   U124 : INVX1 port map( A => Y1(7), Y => n195_port);
   U125 : AND2X1 port map( A => n28, B => 
                           sub_1_root_sub_0_root_sub_184_carry_7_port, Y => 
                           N198);
   U126 : XOR2X1 port map( A => sub_1_root_sub_0_root_sub_184_carry_7_port, B 
                           => n28, Y => N197);
   U127 : AND2X1 port map( A => n29, B => 
                           sub_1_root_sub_0_root_sub_184_carry_6_port, Y => 
                           sub_1_root_sub_0_root_sub_184_carry_7_port);
   U128 : XOR2X1 port map( A => sub_1_root_sub_0_root_sub_184_carry_6_port, B 
                           => n29, Y => N196);
   U129 : AND2X1 port map( A => n30, B => 
                           sub_1_root_sub_0_root_sub_184_carry_5_port, Y => 
                           sub_1_root_sub_0_root_sub_184_carry_6_port);
   U130 : XOR2X1 port map( A => sub_1_root_sub_0_root_sub_184_carry_5_port, B 
                           => n30, Y => N195);
   U131 : AND2X1 port map( A => n31, B => 
                           sub_1_root_sub_0_root_sub_184_carry_4_port, Y => 
                           sub_1_root_sub_0_root_sub_184_carry_5_port);
   U132 : XOR2X1 port map( A => sub_1_root_sub_0_root_sub_184_carry_4_port, B 
                           => n31, Y => N194);
   U133 : AND2X1 port map( A => n32, B => 
                           sub_1_root_sub_0_root_sub_184_carry_3_port, Y => 
                           sub_1_root_sub_0_root_sub_184_carry_4_port);
   U134 : XOR2X1 port map( A => sub_1_root_sub_0_root_sub_184_carry_3_port, B 
                           => n32, Y => N193);
   U135 : AND2X1 port map( A => n33, B => 
                           sub_1_root_sub_0_root_sub_184_carry_2_port, Y => 
                           sub_1_root_sub_0_root_sub_184_carry_3_port);
   U136 : XOR2X1 port map( A => sub_1_root_sub_0_root_sub_184_carry_2_port, B 
                           => n33, Y => N192);
   U137 : AND2X1 port map( A => n34, B => n20, Y => 
                           sub_1_root_sub_0_root_sub_184_carry_2_port);
   U138 : XOR2X1 port map( A => n20, B => n34, Y => N191);
   U139 : INVX2 port map( A => dx_8_port, Y => n28);
   U140 : INVX2 port map( A => n10, Y => n29);
   U141 : INVX2 port map( A => n11, Y => n30);
   U142 : INVX2 port map( A => n12, Y => n31);
   U143 : INVX2 port map( A => n15, Y => n32);
   U144 : INVX2 port map( A => n18, Y => n33);
   U145 : INVX2 port map( A => n19, Y => n34);
   U146 : NAND2X1 port map( A => n44, B => N289, Y => n35);
   U147 : OAI21X1 port map( A => N289, B => n44, C => n35, Y => N290);
   U148 : NOR2X1 port map( A => n35, B => N215, Y => n37);
   U149 : AOI21X1 port map( A => n35, B => N215, C => n37, Y => n36);
   U150 : NAND2X1 port map( A => n37, B => n43, Y => n38);
   U151 : OAI21X1 port map( A => n37, B => n43, C => n38, Y => N292);
   U152 : NOR2X1 port map( A => n38, B => N217, Y => n40);
   U153 : AOI21X1 port map( A => n38, B => N217, C => n40, Y => n39);
   U154 : NAND2X1 port map( A => n40, B => n45, Y => n41);
   U155 : OAI21X1 port map( A => n40, B => n45, C => n41, Y => N294);
   U156 : XNOR2X1 port map( A => N219, B => n41, Y => N295);
   U157 : NOR2X1 port map( A => N219, B => n41, Y => n42);
   U158 : XOR2X1 port map( A => N220, B => n42, Y => N296);
   U159 : INVX2 port map( A => N216, Y => n43);
   U160 : INVX2 port map( A => N214, Y => n44);
   U161 : INVX2 port map( A => N218, Y => n45);
   U162 : INVX2 port map( A => N213, Y => N289);
   U163 : INVX2 port map( A => n39, Y => N293);
   U164 : INVX2 port map( A => n36, Y => N291);
   U165 : NAND2X1 port map( A => n55, B => N326, Y => n46);
   U166 : OAI21X1 port map( A => N326, B => n55, C => n46, Y => N327);
   U167 : NOR2X1 port map( A => n46, B => N231, Y => n48);
   U168 : AOI21X1 port map( A => n46, B => N231, C => n48, Y => n47);
   U169 : NAND2X1 port map( A => n48, B => n54, Y => n49);
   U170 : OAI21X1 port map( A => n48, B => n54, C => n49, Y => N329);
   U171 : NOR2X1 port map( A => n49, B => N209, Y => n51);
   U172 : AOI21X1 port map( A => n49, B => N209, C => n51, Y => n50);
   U173 : NAND2X1 port map( A => n51, B => n56, Y => n52);
   U174 : OAI21X1 port map( A => n51, B => n56, C => n52, Y => N331);
   U175 : XNOR2X1 port map( A => N211, B => n52, Y => N332);
   U176 : NOR2X1 port map( A => N211, B => n52, Y => n53);
   U177 : XOR2X1 port map( A => N212, B => n53, Y => N333);
   U178 : INVX2 port map( A => N232, Y => n54);
   U179 : INVX2 port map( A => N230, Y => n55);
   U180 : INVX2 port map( A => N210, Y => n56);
   U181 : INVX2 port map( A => N229, Y => N326);
   U182 : INVX2 port map( A => n50, Y => N330);
   U183 : INVX2 port map( A => n47, Y => N328);
   U184 : NAND2X1 port map( A => X0(0), B => n152, Y => n58);
   U185 : OAI21X1 port map( A => n58, B => X1(1), C => n153, Y => n57);
   U186 : AOI21X1 port map( A => X1(1), B => n58, C => n154, Y => n59);
   U187 : OAI21X1 port map( A => X0(2), B => n156, C => n59, Y => n60);
   U262 : OAI21X1 port map( A => X1(2), B => n155, C => n60, Y => n61);
   U322 : AOI21X1 port map( A => X0(3), B => n158, C => n61, Y => n62);
   U325 : AOI21X1 port map( A => X1(3), B => n157, C => n62, Y => n63);
   U335 : OAI21X1 port map( A => X0(4), B => n160, C => n63, Y => n64);
   U341 : OAI21X1 port map( A => X1(4), B => n159, C => n64, Y => n65);
   U346 : AOI21X1 port map( A => X0(5), B => n162, C => n65, Y => n66);
   U351 : AOI21X1 port map( A => X1(5), B => n161, C => n66, Y => n67);
   U356 : OAI21X1 port map( A => X0(6), B => n164, C => n67, Y => n149);
   U361 : OAI21X1 port map( A => X1(6), B => n163, C => n149, Y => n150);
   U366 : OAI21X1 port map( A => X0(7), B => n166, C => n150, Y => n151);
   U371 : OAI21X1 port map( A => X1(7), B => n165, C => n151, Y => N95);
   U374 : INVX2 port map( A => X1(0), Y => n152);
   U377 : INVX2 port map( A => X0(1), Y => n153);
   U379 : INVX2 port map( A => n57, Y => n154);
   U381 : INVX2 port map( A => X0(2), Y => n155);
   U387 : INVX2 port map( A => X1(2), Y => n156);
   U392 : INVX2 port map( A => X0(3), Y => n157);
   U397 : INVX2 port map( A => X1(3), Y => n158);
   U402 : INVX2 port map( A => X0(4), Y => n159);
   U407 : INVX2 port map( A => X1(4), Y => n160);
   U412 : INVX2 port map( A => X0(5), Y => n161);
   U417 : INVX2 port map( A => X1(5), Y => n162);
   U420 : INVX2 port map( A => X0(6), Y => n163);
   U421 : INVX2 port map( A => X1(6), Y => n164);
   U427 : INVX2 port map( A => X0(7), Y => n165);
   U429 : INVX2 port map( A => X1(7), Y => n166);
   U514 : NAND2X1 port map( A => Y0(0), B => n181, Y => n168);
   U515 : OAI21X1 port map( A => n168, B => Y1(1), C => n182, Y => n167);
   U516 : AOI21X1 port map( A => Y1(1), B => n168, C => n183, Y => n169);
   U517 : OAI21X1 port map( A => Y0(2), B => n185, C => n169, Y => n170);
   U518 : OAI21X1 port map( A => Y1(2), B => n184, C => n170, Y => n171);
   U519 : AOI21X1 port map( A => Y0(3), B => n187, C => n171, Y => n172);
   U520 : AOI21X1 port map( A => Y1(3), B => n186, C => n172, Y => n173);
   U521 : OAI21X1 port map( A => Y0(4), B => n189, C => n173, Y => n174);
   U522 : OAI21X1 port map( A => Y1(4), B => n188_port, C => n174, Y => n175);
   U523 : AOI21X1 port map( A => Y0(5), B => n191_port, C => n175, Y => n176);
   U524 : AOI21X1 port map( A => Y1(5), B => n190_port, C => n176, Y => n177);
   U525 : OAI21X1 port map( A => Y0(6), B => n193_port, C => n177, Y => n178);
   U526 : OAI21X1 port map( A => Y1(6), B => n192_port, C => n178, Y => n179);
   U527 : OAI21X1 port map( A => Y0(7), B => n195_port, C => n179, Y => n180);
   U528 : OAI21X1 port map( A => Y1(7), B => n194_port, C => n180, Y => N121);
   U529 : INVX2 port map( A => Y1(0), Y => n181);
   U530 : INVX2 port map( A => Y0(1), Y => n182);
   U531 : INVX2 port map( A => n167, Y => n183);
   U532 : INVX2 port map( A => Y0(2), Y => n184);
   U533 : INVX2 port map( A => Y1(2), Y => n185);
   U534 : INVX2 port map( A => Y0(3), Y => n186);
   U535 : INVX2 port map( A => Y1(3), Y => n187);
   U536 : INVX2 port map( A => Y0(4), Y => n188_port);
   U537 : INVX2 port map( A => Y1(4), Y => n189);
   U538 : INVX2 port map( A => Y0(5), Y => n190_port);
   U539 : INVX2 port map( A => Y1(5), Y => n191_port);
   U540 : INVX2 port map( A => Y0(6), Y => n192_port);
   U541 : INVX2 port map( A => Y1(6), Y => n193_port);
   U542 : INVX2 port map( A => Y0(7), Y => n194_port);
   U543 : NAND2X1 port map( A => dy_0_port, B => n220_port, Y => n197_port);
   U544 : OAI21X1 port map( A => n197_port, B => N190, C => n217_port, Y => 
                           n196_port);
   U545 : AOI21X1 port map( A => N190, B => n197_port, C => n221, Y => 
                           n198_port);
   U546 : OAI21X1 port map( A => dy_2_port, B => n34, C => n198_port, Y => 
                           n199_port);
   U547 : OAI21X1 port map( A => n19, B => n216_port, C => n199_port, Y => 
                           n200_port);
   U548 : AOI21X1 port map( A => dy_3_port, B => n33, C => n200_port, Y => 
                           n201_port);
   U549 : AOI21X1 port map( A => n18, B => n215_port, C => n201_port, Y => 
                           n202_port);
   U550 : OAI21X1 port map( A => dy_4_port, B => n32, C => n202_port, Y => 
                           n203_port);
   U551 : OAI21X1 port map( A => n15, B => n214_port, C => n203_port, Y => 
                           n204_port);
   U552 : AOI21X1 port map( A => dy_5_port, B => n31, C => n204_port, Y => 
                           n205_port);
   U553 : AOI21X1 port map( A => n12, B => n213_port, C => n205_port, Y => 
                           n206_port);
   U554 : OAI21X1 port map( A => dy_6_port, B => n30, C => n206_port, Y => 
                           n207_port);
   U555 : OAI21X1 port map( A => n11, B => n212_port, C => n207_port, Y => n208
                           );
   U556 : AOI21X1 port map( A => dy_7_port, B => n29, C => n208, Y => n209_port
                           );
   U557 : AOI21X1 port map( A => n10, B => n218_port, C => n209_port, Y => 
                           n210_port);
   U558 : OAI21X1 port map( A => dy_8_port, B => n28, C => n210_port, Y => 
                           n211_port);
   U559 : OAI21X1 port map( A => dx_8_port, B => n219_port, C => n211_port, Y 
                           => N188);
   U560 : INVX2 port map( A => dy_6_port, Y => n212_port);
   U561 : INVX2 port map( A => dy_5_port, Y => n213_port);
   U562 : INVX2 port map( A => dy_4_port, Y => n214_port);
   U563 : INVX2 port map( A => dy_3_port, Y => n215_port);
   U564 : INVX2 port map( A => dy_2_port, Y => n216_port);
   U565 : INVX2 port map( A => dy_1_port, Y => n217_port);
   U566 : INVX2 port map( A => dy_7_port, Y => n218_port);
   U567 : INVX2 port map( A => dy_8_port, Y => n219_port);
   U568 : INVX2 port map( A => dx_0_port, Y => n220_port);
   U569 : INVX2 port map( A => n196_port, Y => n221);
   U570 : AOI21X1 port map( A => i_1_port, B => n34, C => i_0_port, Y => n222);
   U571 : AOI22X1 port map( A => n222, B => N190, C => n19, D => n561, Y => 
                           n223);
   U572 : OAI21X1 port map( A => i_2_port, B => n33, C => n223, Y => n224);
   U573 : OAI21X1 port map( A => n18, B => n560, C => n224, Y => n225);
   U574 : AOI21X1 port map( A => i_3_port, B => n32, C => n225, Y => n226);
   U575 : AOI21X1 port map( A => n15, B => n559, C => n226, Y => n227);
   U576 : OAI21X1 port map( A => i_4_port, B => n31, C => n227, Y => n228);
   U577 : OAI21X1 port map( A => n12, B => n558, C => n228, Y => n264_port);
   U578 : AOI21X1 port map( A => i_5_port, B => n30, C => n264_port, Y => 
                           n265_port);
   U579 : AOI21X1 port map( A => n11, B => n557, C => n265_port, Y => n361);
   U580 : OAI21X1 port map( A => i_6_port, B => n29, C => n361, Y => n362);
   U581 : OAI21X1 port map( A => n10, B => n556, C => n362, Y => n398);
   U582 : OAI21X1 port map( A => i_7_port, B => n28, C => n398, Y => n399);
   U583 : OAI21X1 port map( A => dx_8_port, B => n562, C => n399, Y => N265);
   U584 : INVX2 port map( A => i_6_port, Y => n556);
   U585 : INVX2 port map( A => i_5_port, Y => n557);
   U586 : INVX2 port map( A => i_4_port, Y => n558);
   U587 : INVX2 port map( A => i_3_port, Y => n559);
   U588 : INVX2 port map( A => i_2_port, Y => n560);
   U589 : INVX2 port map( A => i_1_port, Y => n561);
   U590 : INVX2 port map( A => i_7_port, Y => n562);
   U591 : NOR2X1 port map( A => err_11_port, B => err_10_port, Y => n564);
   U592 : NOR2X1 port map( A => err_9_port, B => err_8_port, Y => n563);
   U593 : NAND2X1 port map( A => n564, B => n563, Y => N266);
   U594 : INVX2 port map( A => N121, Y => n565);
   U595 : INVX2 port map( A => N95, Y => n566);
   U596 : INVX2 port map( A => n476, Y => n567);
   U597 : INVX2 port map( A => n351, Y => n568);
   U598 : INVX2 port map( A => n353, Y => n569);
   U599 : INVX2 port map( A => n354, Y => n570);
   U600 : INVX2 port map( A => n355, Y => n571);
   U601 : INVX2 port map( A => n356, Y => n572);
   U602 : INVX2 port map( A => n357, Y => n573);
   U603 : INVX2 port map( A => n358, Y => n574);
   U604 : INVX2 port map( A => n456, Y => n575);
   U605 : INVX2 port map( A => n479, Y => n577);
   U606 : INVX2 port map( A => n432, Y => n579);
   U607 : INVX2 port map( A => n428, Y => n580);
   U608 : INVX2 port map( A => n424, Y => n581);
   U609 : INVX2 port map( A => n420, Y => n582);
   U610 : INVX2 port map( A => n416, Y => n583);
   U611 : INVX2 port map( A => n412, Y => n584);
   U612 : INVX2 port map( A => n408, Y => n585);
   U613 : INVX2 port map( A => n403, Y => n586);
   U614 : INVX2 port map( A => n392, Y => n587);
   U615 : INVX2 port map( A => n388, Y => n588);
   U616 : INVX2 port map( A => n384, Y => n589);
   U617 : INVX2 port map( A => n380, Y => n590);
   U618 : INVX2 port map( A => n376, Y => n591);
   U619 : INVX2 port map( A => n372, Y => n592);
   U620 : INVX2 port map( A => n367, Y => n593);
   U621 : INVX2 port map( A => n350, Y => n594);
   U622 : INVX2 port map( A => n435, Y => n595);
   U623 : INVX2 port map( A => n480, Y => n596);
   U624 : INVX2 port map( A => n247, Y => rast_done_port);
   U625 : INVX2 port map( A => n245, Y => n598);
   U626 : INVX2 port map( A => n244, Y => n599);
   U627 : INVX2 port map( A => n462, Y => n600);
   U628 : INVX2 port map( A => n436, Y => n602);
   U629 : INVX2 port map( A => state_2_port, Y => n604);
   U630 : INVX2 port map( A => n255, Y => n605);
   U631 : INVX2 port map( A => n298, Y => n608);
   U632 : INVX2 port map( A => n234, Y => n609);
   U633 : INVX2 port map( A => n254, Y => n610);
   U634 : INVX2 port map( A => N188, Y => n613);
   U635 : INVX2 port map( A => err_11_port, Y => n614);
   U636 : INVX2 port map( A => err_10_port, Y => n615);
   U637 : INVX2 port map( A => state_0_port, Y => n616);
   U638 : INVX2 port map( A => n236, Y => n617);
   U639 : INVX2 port map( A => count_3_port, Y => n618);
   U640 : INVX2 port map( A => state_3_port, Y => n619);
   U641 : INVX2 port map( A => n461, Y => n620);
   U642 : INVX2 port map( A => count_0_port, Y => n621);
   U643 : INVX2 port map( A => count_1_port, Y => n622);
   U644 : INVX2 port map( A => count_2_port, Y => n623);
   U645 : INVX2 port map( A => iX, Y => n624);
   U646 : INVX2 port map( A => iY, Y => n625);
   U647 : INVX2 port map( A => err_9_port, Y => n626);
   U648 : INVX2 port map( A => rast_index_1_port, Y => n627);
   U649 : INVX2 port map( A => rast_index_2_port, Y => n628);
   U650 : INVX2 port map( A => rast_index_3_port, Y => n629);
   U651 : INVX2 port map( A => rast_addr_0_port, Y => n630);
   U652 : INVX2 port map( A => rast_addr_1_port, Y => n631);
   U653 : INVX2 port map( A => rast_addr_2_port, Y => n632);
   U654 : INVX2 port map( A => rast_addr_3_port, Y => n633);
   U655 : INVX2 port map( A => rast_addr_4_port, Y => n634);
   U656 : INVX2 port map( A => rast_addr_5_port, Y => n635);
   U657 : INVX2 port map( A => rast_addr_6_port, Y => n636);
   U658 : INVX2 port map( A => rast_addr_7_port, Y => n637);
   U659 : INVX2 port map( A => rast_addr_8_port, Y => n638);
   U660 : INVX2 port map( A => rast_addr_9_port, Y => n639);
   U661 : INVX2 port map( A => rast_addr_10_port, Y => n640);
   U662 : INVX2 port map( A => rast_addr_11_port, Y => n641);
   U663 : INVX2 port map( A => rast_index_0_port, Y => n642);
   U664 : OAI21X1 port map( A => n243, B => n624, C => n255, Y => n349);
   U665 : OAI21X1 port map( A => n243, B => n625, C => n255, Y => n346);
   U666 : NAND2X1 port map( A => N137, B => n404, Y => n405);
   U667 : NAND2X1 port map( A => N136, B => n404, Y => n409);
   U668 : NAND2X1 port map( A => N135, B => n404, Y => n413);
   U669 : NAND2X1 port map( A => N134, B => n404, Y => n417);
   U670 : NAND2X1 port map( A => N133, B => n404, Y => n421);
   U671 : NAND2X1 port map( A => N132, B => n404, Y => n425);
   U672 : NAND2X1 port map( A => N131, B => n404, Y => n429);
   U673 : NAND2X1 port map( A => N138, B => n404, Y => n400);
   U674 : NAND2X1 port map( A => dy_7_port, B => n607, Y => n397);
   U675 : NAND2X1 port map( A => n10, B => n607, Y => n360);
   U676 : NAND2X1 port map( A => N112, B => n368, Y => n364);
   U677 : NAND2X1 port map( A => N111, B => n368, Y => n369);
   U678 : NAND2X1 port map( A => N110, B => n368, Y => n373);
   U679 : NAND2X1 port map( A => N109, B => n368, Y => n377);
   U680 : NAND2X1 port map( A => N108, B => n368, Y => n381);
   U681 : NAND2X1 port map( A => N107, B => n368, Y => n385);
   U682 : NAND2X1 port map( A => N106, B => n368, Y => n389);
   U683 : NAND2X1 port map( A => n255, B => n579, Y => n363);
   U684 : NAND2X1 port map( A => N105, B => n368, Y => n393);
   n643 <= '0';

end SYN_Mixed;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity matrix_math is

   port( screen_cor : out std_logic_vector (7 downto 0);  init_matrix, clk, 
         rst_n : in std_logic;  row_sel : out std_logic_vector (1 downto 0);  
         sel, math_done, strb_screen : out std_logic;  point : in 
         std_logic_vector (47 downto 0);  row : in std_logic_vector (63 downto 
         0);  err : out std_logic);

end matrix_math;

architecture SYN_math_behav of matrix_math is

   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OR2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX2X1
      port( B, A, S : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component BUFX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component matrix_math_DW01_add_18
      port( A, B : in std_logic_vector (23 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (23 downto 0);  CO : out std_logic);
   end component;
   
   component matrix_math_DW01_add_12
      port( A, B : in std_logic_vector (23 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (23 downto 0);  CO : out std_logic);
   end component;
   
   component matrix_math_DW01_add_13
      port( A, B : in std_logic_vector (23 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (23 downto 0);  CO : out std_logic);
   end component;
   
   component matrix_math_DW02_mult_0
      port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (31 downto 0));
   end component;
   
   component matrix_math_DW02_mult_1
      port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (31 downto 0));
   end component;
   
   component matrix_math_DW02_mult_2
      port( A, B : in std_logic_vector (15 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (31 downto 0));
   end component;
   
   component DFFSR
      port( D, CLK, R, S : in std_logic;  Q : out std_logic);
   end component;
   
   signal row_sel_0_port, state_3_port, state_2_port, state_1_port, 
      state_0_port, V1_23_port, n1, n2, n3, n4, n32, n33, n34, n35, N99, N98, 
      N97, N96, N95, N94, N93, N92, N91, N90, N9, N89, N88, N87, N86, N85, N84,
      N83, N82, N81, N80, N8, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70,
      N7, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N6, N59, N58, N57, 
      N56, N55, N54, N53, N52, N51, N50, N5, N49, N48, N47, N46, N45, N44, N43,
      N42, N41, N40, N4_port, N39, N38, N37, N36, N35_port, N34_port, N33_port,
      N32_port, N31, N30, N3_port, N29, N28, N27, N26, N25, N24, N23, N22, N21,
      N20, N2_port, N19, N18, N17, N16, N15, N14, N13, N12, N119, N118, N117, 
      N116, N115, N114, N113, N112, N111, N110, N11, N109, N108, N107, N106, 
      N105, N104, N103, N102, N101, N100, N10, N1_port, N0, n5_port, n6_port, 
      n7_port, n8_port, n9_port, n10_port, n11_port, n12_port, n13_port, 
      n14_port, n15_port, n16_port, n17_port, n18_port, n20_port, n21_port, 
      n22_port, n23_port, n24_port, n25_port, n26_port, n27_port, n28_port, 
      n29_port, n30_port, n31_port, n36_port, n37_port, n38_port, n39_port, 
      n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, 
      n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, 
      n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, 
      n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, 
      n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, 
      n_1273 : std_logic;

begin
   row_sel <= ( n56_port, row_sel_0_port );
   err <= n56_port;
   
   n56_port <= '0';
   state_reg_0_inst : DFFSR port map( D => n48_port, CLK => clk, R => rst_n, S 
                           => n4, Q => state_0_port);
   state_reg_1_inst : DFFSR port map( D => n34, CLK => clk, R => rst_n, S => n3
                           , Q => state_1_port);
   state_reg_2_inst : DFFSR port map( D => n33, CLK => clk, R => rst_n, S => n2
                           , Q => state_2_port);
   state_reg_3_inst : DFFSR port map( D => n14_port, CLK => clk, R => rst_n, S 
                           => n1, Q => state_3_port);
   n1 <= '1';
   n2 <= '1';
   n3 <= '1';
   n4 <= '1';
   U39 : NAND2X1 port map( A => n18_port, B => n12_port, Y => n32);
   mult_53 : matrix_math_DW02_mult_2 port map( A(15) => row(63), A(14) => 
                           row(62), A(13) => row(61), A(12) => row(60), A(11) 
                           => row(59), A(10) => row(58), A(9) => row(57), A(8) 
                           => row(56), A(7) => row(55), A(6) => row(54), A(5) 
                           => row(53), A(4) => row(52), A(3) => row(51), A(2) 
                           => row(50), A(1) => row(49), A(0) => row(48), B(15) 
                           => point(47), B(14) => point(46), B(13) => point(45)
                           , B(12) => point(44), B(11) => point(43), B(10) => 
                           point(42), B(9) => point(41), B(8) => point(40), 
                           B(7) => point(39), B(6) => point(38), B(5) => 
                           point(37), B(4) => point(36), B(3) => point(35), 
                           B(2) => point(34), B(1) => point(33), B(0) => 
                           point(32), TC => n50_port, PRODUCT(31) => n_1231, 
                           PRODUCT(30) => n_1232, PRODUCT(29) => n_1233, 
                           PRODUCT(28) => n_1234, PRODUCT(27) => n_1235, 
                           PRODUCT(26) => n_1236, PRODUCT(25) => n_1237, 
                           PRODUCT(24) => n_1238, PRODUCT(23) => N23, 
                           PRODUCT(22) => N22, PRODUCT(21) => N21, PRODUCT(20) 
                           => N20, PRODUCT(19) => N19, PRODUCT(18) => N18, 
                           PRODUCT(17) => N17, PRODUCT(16) => N16, PRODUCT(15) 
                           => N15, PRODUCT(14) => N14, PRODUCT(13) => N13, 
                           PRODUCT(12) => N12, PRODUCT(11) => N11, PRODUCT(10) 
                           => N10, PRODUCT(9) => N9, PRODUCT(8) => N8, 
                           PRODUCT(7) => N7, PRODUCT(6) => N6, PRODUCT(5) => N5
                           , PRODUCT(4) => N4_port, PRODUCT(3) => N3_port, 
                           PRODUCT(2) => N2_port, PRODUCT(1) => N1_port, 
                           PRODUCT(0) => N0);
   mult_53_2 : matrix_math_DW02_mult_1 port map( A(15) => row(47), A(14) => 
                           row(46), A(13) => row(45), A(12) => row(44), A(11) 
                           => row(43), A(10) => row(42), A(9) => row(41), A(8) 
                           => row(40), A(7) => row(39), A(6) => row(38), A(5) 
                           => row(37), A(4) => row(36), A(3) => row(35), A(2) 
                           => row(34), A(1) => row(33), A(0) => row(32), B(15) 
                           => point(31), B(14) => point(30), B(13) => point(29)
                           , B(12) => point(28), B(11) => point(27), B(10) => 
                           point(26), B(9) => point(25), B(8) => point(24), 
                           B(7) => point(23), B(6) => point(22), B(5) => 
                           point(21), B(4) => point(20), B(3) => point(19), 
                           B(2) => point(18), B(1) => point(17), B(0) => 
                           point(16), TC => n51_port, PRODUCT(31) => n_1239, 
                           PRODUCT(30) => n_1240, PRODUCT(29) => n_1241, 
                           PRODUCT(28) => n_1242, PRODUCT(27) => n_1243, 
                           PRODUCT(26) => n_1244, PRODUCT(25) => n_1245, 
                           PRODUCT(24) => n_1246, PRODUCT(23) => N47, 
                           PRODUCT(22) => N46, PRODUCT(21) => N45, PRODUCT(20) 
                           => N44, PRODUCT(19) => N43, PRODUCT(18) => N42, 
                           PRODUCT(17) => N41, PRODUCT(16) => N40, PRODUCT(15) 
                           => N39, PRODUCT(14) => N38, PRODUCT(13) => N37, 
                           PRODUCT(12) => N36, PRODUCT(11) => N35_port, 
                           PRODUCT(10) => N34_port, PRODUCT(9) => N33_port, 
                           PRODUCT(8) => N32_port, PRODUCT(7) => N31, 
                           PRODUCT(6) => N30, PRODUCT(5) => N29, PRODUCT(4) => 
                           N28, PRODUCT(3) => N27, PRODUCT(2) => N26, 
                           PRODUCT(1) => N25, PRODUCT(0) => N24);
   mult_53_3 : matrix_math_DW02_mult_0 port map( A(15) => row(31), A(14) => 
                           row(30), A(13) => row(29), A(12) => row(28), A(11) 
                           => row(27), A(10) => row(26), A(9) => row(25), A(8) 
                           => row(24), A(7) => row(23), A(6) => row(22), A(5) 
                           => row(21), A(4) => row(20), A(3) => row(19), A(2) 
                           => row(18), A(1) => row(17), A(0) => row(16), B(15) 
                           => point(15), B(14) => point(14), B(13) => point(13)
                           , B(12) => point(12), B(11) => point(11), B(10) => 
                           point(10), B(9) => point(9), B(8) => point(8), B(7) 
                           => point(7), B(6) => point(6), B(5) => point(5), 
                           B(4) => point(4), B(3) => point(3), B(2) => point(2)
                           , B(1) => point(1), B(0) => point(0), TC => n52_port
                           , PRODUCT(31) => n_1247, PRODUCT(30) => n_1248, 
                           PRODUCT(29) => n_1249, PRODUCT(28) => n_1250, 
                           PRODUCT(27) => n_1251, PRODUCT(26) => n_1252, 
                           PRODUCT(25) => n_1253, PRODUCT(24) => n_1254, 
                           PRODUCT(23) => N95, PRODUCT(22) => N94, PRODUCT(21) 
                           => N93, PRODUCT(20) => N92, PRODUCT(19) => N91, 
                           PRODUCT(18) => N90, PRODUCT(17) => N89, PRODUCT(16) 
                           => N88, PRODUCT(15) => N87, PRODUCT(14) => N86, 
                           PRODUCT(13) => N85, PRODUCT(12) => N84, PRODUCT(11) 
                           => N83, PRODUCT(10) => N82, PRODUCT(9) => N81, 
                           PRODUCT(8) => N80, PRODUCT(7) => N79, PRODUCT(6) => 
                           N78, PRODUCT(5) => N77, PRODUCT(4) => N76, 
                           PRODUCT(3) => N75, PRODUCT(2) => N74, PRODUCT(1) => 
                           N73, PRODUCT(0) => N72);
   add_1_root_add_0_root_add_53_3 : matrix_math_DW01_add_13 port map( A(23) => 
                           N23, A(22) => N22, A(21) => N21, A(20) => N20, A(19)
                           => N19, A(18) => N18, A(17) => N17, A(16) => N16, 
                           A(15) => N15, A(14) => N14, A(13) => N13, A(12) => 
                           N12, A(11) => N11, A(10) => N10, A(9) => N9, A(8) =>
                           N8, A(7) => N7, A(6) => N6, A(5) => N5, A(4) => 
                           N4_port, A(3) => N3_port, A(2) => N2_port, A(1) => 
                           N1_port, A(0) => N0, B(23) => N95, B(22) => N94, 
                           B(21) => N93, B(20) => N92, B(19) => N91, B(18) => 
                           N90, B(17) => N89, B(16) => N88, B(15) => N87, B(14)
                           => N86, B(13) => N85, B(12) => N84, B(11) => N83, 
                           B(10) => N82, B(9) => N81, B(8) => N80, B(7) => N79,
                           B(6) => N78, B(5) => N77, B(4) => N76, B(3) => N75, 
                           B(2) => N74, B(1) => N73, B(0) => N72, CI => 
                           n53_port, SUM(23) => N71, SUM(22) => N70, SUM(21) =>
                           N69, SUM(20) => N68, SUM(19) => N67, SUM(18) => N66,
                           SUM(17) => N65, SUM(16) => N64, SUM(15) => N63, 
                           SUM(14) => N62, SUM(13) => N61, SUM(12) => N60, 
                           SUM(11) => N59, SUM(10) => N58, SUM(9) => N57, 
                           SUM(8) => N56, SUM(7) => N55, SUM(6) => N54, SUM(5) 
                           => N53, SUM(4) => N52, SUM(3) => N51, SUM(2) => N50,
                           SUM(1) => N49, SUM(0) => N48, CO => n_1255);
   add_2_root_add_0_root_add_53_3 : matrix_math_DW01_add_12 port map( A(23) => 
                           row(15), A(22) => row(14), A(21) => row(13), A(20) 
                           => row(12), A(19) => row(11), A(18) => row(10), 
                           A(17) => row(9), A(16) => row(8), A(15) => row(7), 
                           A(14) => row(6), A(13) => row(5), A(12) => row(4), 
                           A(11) => row(3), A(10) => row(2), A(9) => row(1), 
                           A(8) => row(0), A(7) => n49_port, A(6) => n49_port, 
                           A(5) => n49_port, A(4) => n49_port, A(3) => n49_port
                           , A(2) => n49_port, A(1) => n49_port, A(0) => 
                           n49_port, B(23) => N47, B(22) => N46, B(21) => N45, 
                           B(20) => N44, B(19) => N43, B(18) => N42, B(17) => 
                           N41, B(16) => N40, B(15) => N39, B(14) => N38, B(13)
                           => N37, B(12) => N36, B(11) => N35_port, B(10) => 
                           N34_port, B(9) => N33_port, B(8) => N32_port, B(7) 
                           => N31, B(6) => N30, B(5) => N29, B(4) => N28, B(3) 
                           => N27, B(2) => N26, B(1) => N25, B(0) => N24, CI =>
                           n54_port, SUM(23) => N119, SUM(22) => N118, SUM(21) 
                           => N117, SUM(20) => N116, SUM(19) => N115, SUM(18) 
                           => N114, SUM(17) => N113, SUM(16) => N112, SUM(15) 
                           => N111, SUM(14) => N110, SUM(13) => N109, SUM(12) 
                           => N108, SUM(11) => N107, SUM(10) => N106, SUM(9) =>
                           N105, SUM(8) => N104, SUM(7) => N103, SUM(6) => N102
                           , SUM(5) => N101, SUM(4) => N100, SUM(3) => N99, 
                           SUM(2) => N98, SUM(1) => N97, SUM(0) => N96, CO => 
                           n_1256);
   add_0_root_add_0_root_add_53_3 : matrix_math_DW01_add_18 port map( A(23) => 
                           N71, A(22) => N70, A(21) => N69, A(20) => N68, A(19)
                           => N67, A(18) => N66, A(17) => N65, A(16) => N64, 
                           A(15) => N63, A(14) => N62, A(13) => N61, A(12) => 
                           N60, A(11) => N59, A(10) => N58, A(9) => N57, A(8) 
                           => N56, A(7) => N55, A(6) => N54, A(5) => N53, A(4) 
                           => N52, A(3) => N51, A(2) => N50, A(1) => N49, A(0) 
                           => N48, B(23) => N119, B(22) => N118, B(21) => N117,
                           B(20) => N116, B(19) => N115, B(18) => N114, B(17) 
                           => N113, B(16) => N112, B(15) => N111, B(14) => N110
                           , B(13) => N109, B(12) => N108, B(11) => N107, B(10)
                           => N106, B(9) => N105, B(8) => N104, B(7) => N103, 
                           B(6) => N102, B(5) => N101, B(4) => N100, B(3) => 
                           N99, B(2) => N98, B(1) => N97, B(0) => N96, CI => 
                           n55_port, SUM(23) => V1_23_port, SUM(22) => 
                           screen_cor(6), SUM(21) => screen_cor(5), SUM(20) => 
                           screen_cor(4), SUM(19) => screen_cor(3), SUM(18) => 
                           screen_cor(2), SUM(17) => screen_cor(1), SUM(16) => 
                           screen_cor(0), SUM(15) => n_1257, SUM(14) => n_1258,
                           SUM(13) => n_1259, SUM(12) => n_1260, SUM(11) => 
                           n_1261, SUM(10) => n_1262, SUM(9) => n_1263, SUM(8) 
                           => n_1264, SUM(7) => n_1265, SUM(6) => n_1266, 
                           SUM(5) => n_1267, SUM(4) => n_1268, SUM(3) => n_1269
                           , SUM(2) => n_1270, SUM(1) => n_1271, SUM(0) => 
                           n_1272, CO => n_1273);
   U6 : BUFX2 port map( A => n22_port, Y => n5_port);
   U7 : BUFX2 port map( A => state_1_port, Y => n6_port);
   U8 : INVX1 port map( A => state_1_port, Y => n17_port);
   U9 : BUFX4 port map( A => state_0_port, Y => n7_port);
   U10 : BUFX2 port map( A => state_0_port, Y => n16_port);
   U11 : INVX2 port map( A => n17_port, Y => n8_port);
   U12 : INVX1 port map( A => n28_port, Y => n9_port);
   U13 : INVX1 port map( A => n35, Y => n36_port);
   U14 : INVX2 port map( A => state_2_port, Y => n10_port);
   U15 : INVX4 port map( A => n10_port, Y => n11_port);
   U16 : BUFX4 port map( A => state_3_port, Y => n12_port);
   U17 : INVX1 port map( A => state_3_port, Y => n39_port);
   U18 : BUFX2 port map( A => n8_port, Y => n13_port);
   U19 : OAI21X1 port map( A => n24_port, B => n23_port, C => n22_port, Y => 
                           n14_port);
   U20 : INVX2 port map( A => n15_port, Y => strb_screen);
   U21 : AND2X2 port map( A => n21_port, B => n5_port, Y => n15_port);
   U22 : BUFX2 port map( A => n7_port, Y => n18_port);
   U23 : INVX1 port map( A => n6_port, Y => n24_port);
   U24 : OR2X2 port map( A => n18_port, B => n12_port, Y => n46_port);
   U25 : INVX2 port map( A => n46_port, Y => n41_port);
   U26 : OR2X2 port map( A => n13_port, B => n11_port, Y => n38_port);
   U27 : NAND2X1 port map( A => n41_port, B => n38_port, Y => n21_port);
   U28 : INVX2 port map( A => n11_port, Y => n29_port);
   U29 : NOR2X1 port map( A => n6_port, B => n16_port, Y => n20_port);
   U30 : NAND3X1 port map( A => n12_port, B => n29_port, C => n20_port, Y => 
                           n22_port);
   U31 : NOR2X1 port map( A => n32, B => n38_port, Y => math_done);
   U32 : NAND3X1 port map( A => n11_port, B => n7_port, C => n39_port, Y => 
                           n23_port);
   U33 : OAI21X1 port map( A => n24_port, B => n23_port, C => n22_port, Y => 
                           n35);
   U34 : NAND2X1 port map( A => n6_port, B => n16_port, Y => n25_port);
   U35 : NOR2X1 port map( A => n12_port, B => n25_port, Y => n27_port);
   U36 : NOR3X1 port map( A => n7_port, B => n12_port, C => n8_port, Y => 
                           n26_port);
   U37 : MUX2X1 port map( B => n27_port, A => n26_port, S => n11_port, Y => 
                           n37_port);
   U38 : INVX2 port map( A => n37_port, Y => n28_port);
   U40 : OR2X2 port map( A => n28_port, B => n14_port, Y => sel);
   U41 : NOR2X1 port map( A => n12_port, B => n29_port, Y => n31_port);
   U42 : XOR2X1 port map( A => n7_port, B => n8_port, Y => n30_port);
   U43 : NAND2X1 port map( A => n31_port, B => n30_port, Y => n43_port);
   U44 : NAND2X1 port map( A => n36_port, B => n43_port, Y => row_sel_0_port);
   U45 : INVX2 port map( A => V1_23_port, Y => screen_cor(7));
   U46 : NAND2X1 port map( A => n43_port, B => n9_port, Y => n33);
   U47 : INVX2 port map( A => n38_port, Y => n40_port);
   U48 : NAND3X1 port map( A => n18_port, B => n40_port, C => n39_port, Y => 
                           n44_port);
   U49 : NAND2X1 port map( A => n13_port, B => n41_port, Y => n42_port);
   U50 : NAND3X1 port map( A => n44_port, B => n43_port, C => n42_port, Y => 
                           n34);
   U51 : INVX2 port map( A => init_matrix, Y => n45_port);
   U52 : OAI21X1 port map( A => n46_port, B => n45_port, C => n15_port, Y => 
                           n48_port);
   n49_port <= '0';
   n50_port <= '1';
   n51_port <= '1';
   n52_port <= '1';
   n53_port <= '0';
   n54_port <= '0';
   n55_port <= '0';

end SYN_math_behav;

library IEEE,OSU_AMI05;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_overall.all;

entity overall is

   port( databus : inout std_logic_vector (15 downto 0);  addr_out : out 
         std_logic_vector (14 downto 0);  re_out, we_out : out std_logic;  
         strb_in, ram_in_use : in std_logic;  gpu_done : out std_logic;  clk, 
         rst_n : in std_logic);

end overall;

architecture SYN_struct of overall is

   component gpu_controller
      port( databus : inout std_logic_vector (15 downto 0);  strb_in, clk, 
            rst_n : in std_logic;  gpu_done : out std_logic;  ram_in_use, 
            rast_done : in std_logic;  init_rast : out std_logic;  rast_addr : 
            in std_logic_vector (15 downto 0);  rast_strb : in std_logic;  
            rast_index : in std_logic_vector (3 downto 0);  math_done : in 
            std_logic;  init_math, strb_matrix, strb_cor : out std_logic;  err 
            : in std_logic;  addr_out : out std_logic_vector (14 downto 0);  
            re_out, we_out : out std_logic;  databus_out, opp : out 
            std_logic_vector (15 downto 0));
   end component;
   
   component coordinate_buffer
      port( strb_cor : in std_logic;  databus_out : in std_logic_vector (15 
            downto 0);  clk, sel : in std_logic;  point : out std_logic_vector 
            (47 downto 0));
   end component;
   
   component world_matrix_buffer
      port( strb_matrix : in std_logic;  databus_out : in std_logic_vector (15 
            downto 0);  clk : in std_logic;  row_sel : in std_logic_vector (1 
            downto 0);  row : out std_logic_vector (63 downto 0));
   end component;
   
   component screen_buffer
      port( clk, strb_screen : in std_logic;  screen_cor : in std_logic_vector 
            (7 downto 0);  X0, X1, Y0, Y1 : out std_logic_vector (7 downto 0));
   end component;
   
   component Rasterizer
      port( clk : in std_logic;  X0, X1, Y0, Y1 : in std_logic_vector (7 downto
            0);  init_rast, RST_N : in std_logic;  rast_done, rast_strb : out 
            std_logic;  rast_index : out std_logic_vector (3 downto 0);  
            rast_addr : out std_logic_vector (15 downto 0));
   end component;
   
   component matrix_math
      port( screen_cor : out std_logic_vector (7 downto 0);  init_matrix, clk, 
            rst_n : in std_logic;  row_sel : out std_logic_vector (1 downto 0);
            sel, math_done, strb_screen : out std_logic;  point : in 
            std_logic_vector (47 downto 0);  row : in std_logic_vector (63 
            downto 0);  err : out std_logic);
   end component;
   
   signal math_done, init_math, point_47_port, point_46_port, point_45_port, 
      point_44_port, point_43_port, point_42_port, point_41_port, point_40_port
      , point_39_port, point_38_port, point_37_port, point_36_port, 
      point_35_port, point_34_port, point_33_port, point_32_port, point_31_port
      , point_30_port, point_29_port, point_28_port, point_27_port, 
      point_26_port, point_25_port, point_24_port, point_23_port, point_22_port
      , point_21_port, point_20_port, point_19_port, point_18_port, 
      point_17_port, point_16_port, point_15_port, point_14_port, point_13_port
      , point_12_port, point_11_port, point_10_port, point_9_port, point_8_port
      , point_7_port, point_6_port, point_5_port, point_4_port, point_3_port, 
      point_2_port, point_1_port, point_0_port, row_63_port, row_62_port, 
      row_61_port, row_60_port, row_59_port, row_58_port, row_57_port, 
      row_56_port, row_55_port, row_54_port, row_53_port, row_52_port, 
      row_51_port, row_50_port, row_49_port, row_48_port, row_47_port, 
      row_46_port, row_45_port, row_44_port, row_43_port, row_42_port, 
      row_41_port, row_40_port, row_39_port, row_38_port, row_37_port, 
      row_36_port, row_35_port, row_34_port, row_33_port, row_32_port, 
      row_31_port, row_30_port, row_29_port, row_28_port, row_27_port, 
      row_26_port, row_25_port, row_24_port, row_23_port, row_22_port, 
      row_21_port, row_20_port, row_19_port, row_18_port, row_17_port, 
      row_16_port, row_15_port, row_14_port, row_13_port, row_12_port, 
      row_11_port, row_10_port, row_9_port, row_8_port, row_7_port, row_6_port,
      row_5_port, row_4_port, row_3_port, row_2_port, row_1_port, row_0_port, 
      screen_cor_7_port, screen_cor_6_port, screen_cor_5_port, 
      screen_cor_4_port, screen_cor_3_port, screen_cor_2_port, 
      screen_cor_1_port, screen_cor_0_port, strb_screen, row_sel_1_port, 
      row_sel_0_port, err, sel, X0_7_port, X0_6_port, X0_5_port, X0_4_port, 
      X0_3_port, X0_2_port, X0_1_port, X0_0_port, X1_7_port, X1_6_port, 
      X1_5_port, X1_4_port, X1_3_port, X1_2_port, X1_1_port, X1_0_port, 
      Y0_7_port, Y0_6_port, Y0_5_port, Y0_4_port, Y0_3_port, Y0_2_port, 
      Y0_1_port, Y0_0_port, Y1_7_port, Y1_6_port, Y1_5_port, Y1_4_port, 
      Y1_3_port, Y1_2_port, Y1_1_port, Y1_0_port, init_rast, rast_done, 
      rast_strb, rast_index_3_port, rast_index_2_port, rast_index_1_port, 
      rast_index_0_port, rast_addr_15_port, rast_addr_14_port, 
      rast_addr_13_port, rast_addr_12_port, rast_addr_11_port, 
      rast_addr_10_port, rast_addr_9_port, rast_addr_8_port, rast_addr_7_port, 
      rast_addr_6_port, rast_addr_5_port, rast_addr_4_port, rast_addr_3_port, 
      rast_addr_2_port, rast_addr_1_port, rast_addr_0_port, strb_matrix, 
      databus_out_15_port, databus_out_14_port, databus_out_13_port, 
      databus_out_12_port, databus_out_11_port, databus_out_10_port, 
      databus_out_9_port, databus_out_8_port, databus_out_7_port, 
      databus_out_6_port, databus_out_5_port, databus_out_4_port, 
      databus_out_3_port, databus_out_2_port, databus_out_1_port, 
      databus_out_0_port, strb_cor, n_1274, n_1275, n_1276, n_1277, n_1278, 
      n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, 
      n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295 : 
      std_logic;

begin
   
   DUT5 : matrix_math port map( screen_cor(7) => screen_cor_7_port, 
                           screen_cor(6) => screen_cor_6_port, screen_cor(5) =>
                           screen_cor_5_port, screen_cor(4) => 
                           screen_cor_4_port, screen_cor(3) => 
                           screen_cor_3_port, screen_cor(2) => 
                           screen_cor_2_port, screen_cor(1) => 
                           screen_cor_1_port, screen_cor(0) => 
                           screen_cor_0_port, init_matrix => init_math, clk => 
                           clk, rst_n => rst_n, row_sel(1) => n_1274, 
                           row_sel(0) => row_sel_0_port, sel => sel, math_done 
                           => math_done, strb_screen => strb_screen, point(47) 
                           => point_47_port, point(46) => point_46_port, 
                           point(45) => point_45_port, point(44) => 
                           point_44_port, point(43) => point_43_port, point(42)
                           => point_42_port, point(41) => point_41_port, 
                           point(40) => point_40_port, point(39) => 
                           point_39_port, point(38) => point_38_port, point(37)
                           => point_37_port, point(36) => point_36_port, 
                           point(35) => point_35_port, point(34) => 
                           point_34_port, point(33) => point_33_port, point(32)
                           => point_32_port, point(31) => point_31_port, 
                           point(30) => point_30_port, point(29) => 
                           point_29_port, point(28) => point_28_port, point(27)
                           => point_27_port, point(26) => point_26_port, 
                           point(25) => point_25_port, point(24) => 
                           point_24_port, point(23) => point_23_port, point(22)
                           => point_22_port, point(21) => point_21_port, 
                           point(20) => point_20_port, point(19) => 
                           point_19_port, point(18) => point_18_port, point(17)
                           => point_17_port, point(16) => point_16_port, 
                           point(15) => point_15_port, point(14) => 
                           point_14_port, point(13) => point_13_port, point(12)
                           => point_12_port, point(11) => point_11_port, 
                           point(10) => point_10_port, point(9) => point_9_port
                           , point(8) => point_8_port, point(7) => point_7_port
                           , point(6) => point_6_port, point(5) => point_5_port
                           , point(4) => point_4_port, point(3) => point_3_port
                           , point(2) => point_2_port, point(1) => point_1_port
                           , point(0) => point_0_port, row(63) => row_63_port, 
                           row(62) => row_62_port, row(61) => row_61_port, 
                           row(60) => row_60_port, row(59) => row_59_port, 
                           row(58) => row_58_port, row(57) => row_57_port, 
                           row(56) => row_56_port, row(55) => row_55_port, 
                           row(54) => row_54_port, row(53) => row_53_port, 
                           row(52) => row_52_port, row(51) => row_51_port, 
                           row(50) => row_50_port, row(49) => row_49_port, 
                           row(48) => row_48_port, row(47) => row_47_port, 
                           row(46) => row_46_port, row(45) => row_45_port, 
                           row(44) => row_44_port, row(43) => row_43_port, 
                           row(42) => row_42_port, row(41) => row_41_port, 
                           row(40) => row_40_port, row(39) => row_39_port, 
                           row(38) => row_38_port, row(37) => row_37_port, 
                           row(36) => row_36_port, row(35) => row_35_port, 
                           row(34) => row_34_port, row(33) => row_33_port, 
                           row(32) => row_32_port, row(31) => row_31_port, 
                           row(30) => row_30_port, row(29) => row_29_port, 
                           row(28) => row_28_port, row(27) => row_27_port, 
                           row(26) => row_26_port, row(25) => row_25_port, 
                           row(24) => row_24_port, row(23) => row_23_port, 
                           row(22) => row_22_port, row(21) => row_21_port, 
                           row(20) => row_20_port, row(19) => row_19_port, 
                           row(18) => row_18_port, row(17) => row_17_port, 
                           row(16) => row_16_port, row(15) => row_15_port, 
                           row(14) => row_14_port, row(13) => row_13_port, 
                           row(12) => row_12_port, row(11) => row_11_port, 
                           row(10) => row_10_port, row(9) => row_9_port, row(8)
                           => row_8_port, row(7) => row_7_port, row(6) => 
                           row_6_port, row(5) => row_5_port, row(4) => 
                           row_4_port, row(3) => row_3_port, row(2) => 
                           row_2_port, row(1) => row_1_port, row(0) => 
                           row_0_port, err => n_1275);
   DUT4 : Rasterizer port map( clk => clk, X0(7) => X0_7_port, X0(6) => 
                           X0_6_port, X0(5) => X0_5_port, X0(4) => X0_4_port, 
                           X0(3) => X0_3_port, X0(2) => X0_2_port, X0(1) => 
                           X0_1_port, X0(0) => X0_0_port, X1(7) => X1_7_port, 
                           X1(6) => X1_6_port, X1(5) => X1_5_port, X1(4) => 
                           X1_4_port, X1(3) => X1_3_port, X1(2) => X1_2_port, 
                           X1(1) => X1_1_port, X1(0) => X1_0_port, Y0(7) => 
                           Y0_7_port, Y0(6) => Y0_6_port, Y0(5) => Y0_5_port, 
                           Y0(4) => Y0_4_port, Y0(3) => Y0_3_port, Y0(2) => 
                           Y0_2_port, Y0(1) => Y0_1_port, Y0(0) => Y0_0_port, 
                           Y1(7) => Y1_7_port, Y1(6) => Y1_6_port, Y1(5) => 
                           Y1_5_port, Y1(4) => Y1_4_port, Y1(3) => Y1_3_port, 
                           Y1(2) => Y1_2_port, Y1(1) => Y1_1_port, Y1(0) => 
                           Y1_0_port, init_rast => init_rast, RST_N => rst_n, 
                           rast_done => rast_done, rast_strb => rast_strb, 
                           rast_index(3) => rast_index_3_port, rast_index(2) =>
                           rast_index_2_port, rast_index(1) => 
                           rast_index_1_port, rast_index(0) => 
                           rast_index_0_port, rast_addr(15) => n_1276, 
                           rast_addr(14) => n_1277, rast_addr(13) => n_1278, 
                           rast_addr(12) => n_1279, rast_addr(11) => 
                           rast_addr_11_port, rast_addr(10) => 
                           rast_addr_10_port, rast_addr(9) => rast_addr_9_port,
                           rast_addr(8) => rast_addr_8_port, rast_addr(7) => 
                           rast_addr_7_port, rast_addr(6) => rast_addr_6_port, 
                           rast_addr(5) => rast_addr_5_port, rast_addr(4) => 
                           rast_addr_4_port, rast_addr(3) => rast_addr_3_port, 
                           rast_addr(2) => rast_addr_2_port, rast_addr(1) => 
                           rast_addr_1_port, rast_addr(0) => rast_addr_0_port);
   DUT3 : screen_buffer port map( clk => clk, strb_screen => strb_screen, 
                           screen_cor(7) => screen_cor_7_port, screen_cor(6) =>
                           screen_cor_6_port, screen_cor(5) => 
                           screen_cor_5_port, screen_cor(4) => 
                           screen_cor_4_port, screen_cor(3) => 
                           screen_cor_3_port, screen_cor(2) => 
                           screen_cor_2_port, screen_cor(1) => 
                           screen_cor_1_port, screen_cor(0) => 
                           screen_cor_0_port, X0(7) => X0_7_port, X0(6) => 
                           X0_6_port, X0(5) => X0_5_port, X0(4) => X0_4_port, 
                           X0(3) => X0_3_port, X0(2) => X0_2_port, X0(1) => 
                           X0_1_port, X0(0) => X0_0_port, X1(7) => X1_7_port, 
                           X1(6) => X1_6_port, X1(5) => X1_5_port, X1(4) => 
                           X1_4_port, X1(3) => X1_3_port, X1(2) => X1_2_port, 
                           X1(1) => X1_1_port, X1(0) => X1_0_port, Y0(7) => 
                           Y0_7_port, Y0(6) => Y0_6_port, Y0(5) => Y0_5_port, 
                           Y0(4) => Y0_4_port, Y0(3) => Y0_3_port, Y0(2) => 
                           Y0_2_port, Y0(1) => Y0_1_port, Y0(0) => Y0_0_port, 
                           Y1(7) => Y1_7_port, Y1(6) => Y1_6_port, Y1(5) => 
                           Y1_5_port, Y1(4) => Y1_4_port, Y1(3) => Y1_3_port, 
                           Y1(2) => Y1_2_port, Y1(1) => Y1_1_port, Y1(0) => 
                           Y1_0_port);
   DUT2 : world_matrix_buffer port map( strb_matrix => strb_matrix, 
                           databus_out(15) => databus_out_15_port, 
                           databus_out(14) => databus_out_14_port, 
                           databus_out(13) => databus_out_13_port, 
                           databus_out(12) => databus_out_12_port, 
                           databus_out(11) => databus_out_11_port, 
                           databus_out(10) => databus_out_10_port, 
                           databus_out(9) => databus_out_9_port, databus_out(8)
                           => databus_out_8_port, databus_out(7) => 
                           databus_out_7_port, databus_out(6) => 
                           databus_out_6_port, databus_out(5) => 
                           databus_out_5_port, databus_out(4) => 
                           databus_out_4_port, databus_out(3) => 
                           databus_out_3_port, databus_out(2) => 
                           databus_out_2_port, databus_out(1) => 
                           databus_out_1_port, databus_out(0) => 
                           databus_out_0_port, clk => clk, row_sel(1) => 
                           row_sel_1_port, row_sel(0) => row_sel_0_port, 
                           row(63) => row_63_port, row(62) => row_62_port, 
                           row(61) => row_61_port, row(60) => row_60_port, 
                           row(59) => row_59_port, row(58) => row_58_port, 
                           row(57) => row_57_port, row(56) => row_56_port, 
                           row(55) => row_55_port, row(54) => row_54_port, 
                           row(53) => row_53_port, row(52) => row_52_port, 
                           row(51) => row_51_port, row(50) => row_50_port, 
                           row(49) => row_49_port, row(48) => row_48_port, 
                           row(47) => row_47_port, row(46) => row_46_port, 
                           row(45) => row_45_port, row(44) => row_44_port, 
                           row(43) => row_43_port, row(42) => row_42_port, 
                           row(41) => row_41_port, row(40) => row_40_port, 
                           row(39) => row_39_port, row(38) => row_38_port, 
                           row(37) => row_37_port, row(36) => row_36_port, 
                           row(35) => row_35_port, row(34) => row_34_port, 
                           row(33) => row_33_port, row(32) => row_32_port, 
                           row(31) => row_31_port, row(30) => row_30_port, 
                           row(29) => row_29_port, row(28) => row_28_port, 
                           row(27) => row_27_port, row(26) => row_26_port, 
                           row(25) => row_25_port, row(24) => row_24_port, 
                           row(23) => row_23_port, row(22) => row_22_port, 
                           row(21) => row_21_port, row(20) => row_20_port, 
                           row(19) => row_19_port, row(18) => row_18_port, 
                           row(17) => row_17_port, row(16) => row_16_port, 
                           row(15) => row_15_port, row(14) => row_14_port, 
                           row(13) => row_13_port, row(12) => row_12_port, 
                           row(11) => row_11_port, row(10) => row_10_port, 
                           row(9) => row_9_port, row(8) => row_8_port, row(7) 
                           => row_7_port, row(6) => row_6_port, row(5) => 
                           row_5_port, row(4) => row_4_port, row(3) => 
                           row_3_port, row(2) => row_2_port, row(1) => 
                           row_1_port, row(0) => row_0_port);
   DUT1 : coordinate_buffer port map( strb_cor => strb_cor, databus_out(15) => 
                           databus_out_15_port, databus_out(14) => 
                           databus_out_14_port, databus_out(13) => 
                           databus_out_13_port, databus_out(12) => 
                           databus_out_12_port, databus_out(11) => 
                           databus_out_11_port, databus_out(10) => 
                           databus_out_10_port, databus_out(9) => 
                           databus_out_9_port, databus_out(8) => 
                           databus_out_8_port, databus_out(7) => 
                           databus_out_7_port, databus_out(6) => 
                           databus_out_6_port, databus_out(5) => 
                           databus_out_5_port, databus_out(4) => 
                           databus_out_4_port, databus_out(3) => 
                           databus_out_3_port, databus_out(2) => 
                           databus_out_2_port, databus_out(1) => 
                           databus_out_1_port, databus_out(0) => 
                           databus_out_0_port, clk => clk, sel => sel, 
                           point(47) => point_47_port, point(46) => 
                           point_46_port, point(45) => point_45_port, point(44)
                           => point_44_port, point(43) => point_43_port, 
                           point(42) => point_42_port, point(41) => 
                           point_41_port, point(40) => point_40_port, point(39)
                           => point_39_port, point(38) => point_38_port, 
                           point(37) => point_37_port, point(36) => 
                           point_36_port, point(35) => point_35_port, point(34)
                           => point_34_port, point(33) => point_33_port, 
                           point(32) => point_32_port, point(31) => 
                           point_31_port, point(30) => point_30_port, point(29)
                           => point_29_port, point(28) => point_28_port, 
                           point(27) => point_27_port, point(26) => 
                           point_26_port, point(25) => point_25_port, point(24)
                           => point_24_port, point(23) => point_23_port, 
                           point(22) => point_22_port, point(21) => 
                           point_21_port, point(20) => point_20_port, point(19)
                           => point_19_port, point(18) => point_18_port, 
                           point(17) => point_17_port, point(16) => 
                           point_16_port, point(15) => point_15_port, point(14)
                           => point_14_port, point(13) => point_13_port, 
                           point(12) => point_12_port, point(11) => 
                           point_11_port, point(10) => point_10_port, point(9) 
                           => point_9_port, point(8) => point_8_port, point(7) 
                           => point_7_port, point(6) => point_6_port, point(5) 
                           => point_5_port, point(4) => point_4_port, point(3) 
                           => point_3_port, point(2) => point_2_port, point(1) 
                           => point_1_port, point(0) => point_0_port);
   DUT : gpu_controller port map( databus(15) => databus(15), databus(14) => 
                           databus(14), databus(13) => databus(13), databus(12)
                           => databus(12), databus(11) => databus(11), 
                           databus(10) => databus(10), databus(9) => databus(9)
                           , databus(8) => databus(8), databus(7) => databus(7)
                           , databus(6) => databus(6), databus(5) => databus(5)
                           , databus(4) => databus(4), databus(3) => databus(3)
                           , databus(2) => databus(2), databus(1) => databus(1)
                           , databus(0) => databus(0), strb_in => strb_in, clk 
                           => clk, rst_n => rst_n, gpu_done => gpu_done, 
                           ram_in_use => ram_in_use, rast_done => rast_done, 
                           init_rast => init_rast, rast_addr(15) => 
                           rast_addr_15_port, rast_addr(14) => 
                           rast_addr_14_port, rast_addr(13) => 
                           rast_addr_13_port, rast_addr(12) => 
                           rast_addr_12_port, rast_addr(11) => 
                           rast_addr_11_port, rast_addr(10) => 
                           rast_addr_10_port, rast_addr(9) => rast_addr_9_port,
                           rast_addr(8) => rast_addr_8_port, rast_addr(7) => 
                           rast_addr_7_port, rast_addr(6) => rast_addr_6_port, 
                           rast_addr(5) => rast_addr_5_port, rast_addr(4) => 
                           rast_addr_4_port, rast_addr(3) => rast_addr_3_port, 
                           rast_addr(2) => rast_addr_2_port, rast_addr(1) => 
                           rast_addr_1_port, rast_addr(0) => rast_addr_0_port, 
                           rast_strb => rast_strb, rast_index(3) => 
                           rast_index_3_port, rast_index(2) => 
                           rast_index_2_port, rast_index(1) => 
                           rast_index_1_port, rast_index(0) => 
                           rast_index_0_port, math_done => math_done, init_math
                           => init_math, strb_matrix => strb_matrix, strb_cor 
                           => strb_cor, err => err, addr_out(14) => 
                           addr_out(14), addr_out(13) => addr_out(13), 
                           addr_out(12) => addr_out(12), addr_out(11) => 
                           addr_out(11), addr_out(10) => addr_out(10), 
                           addr_out(9) => addr_out(9), addr_out(8) => 
                           addr_out(8), addr_out(7) => addr_out(7), addr_out(6)
                           => addr_out(6), addr_out(5) => addr_out(5), 
                           addr_out(4) => addr_out(4), addr_out(3) => 
                           addr_out(3), addr_out(2) => addr_out(2), addr_out(1)
                           => addr_out(1), addr_out(0) => addr_out(0), re_out 
                           => re_out, we_out => we_out, databus_out(15) => 
                           databus_out_15_port, databus_out(14) => 
                           databus_out_14_port, databus_out(13) => 
                           databus_out_13_port, databus_out(12) => 
                           databus_out_12_port, databus_out(11) => 
                           databus_out_11_port, databus_out(10) => 
                           databus_out_10_port, databus_out(9) => 
                           databus_out_9_port, databus_out(8) => 
                           databus_out_8_port, databus_out(7) => 
                           databus_out_7_port, databus_out(6) => 
                           databus_out_6_port, databus_out(5) => 
                           databus_out_5_port, databus_out(4) => 
                           databus_out_4_port, databus_out(3) => 
                           databus_out_3_port, databus_out(2) => 
                           databus_out_2_port, databus_out(1) => 
                           databus_out_1_port, databus_out(0) => 
                           databus_out_0_port, opp(15) => n_1280, opp(14) => 
                           n_1281, opp(13) => n_1282, opp(12) => n_1283, 
                           opp(11) => n_1284, opp(10) => n_1285, opp(9) => 
                           n_1286, opp(8) => n_1287, opp(7) => n_1288, opp(6) 
                           => n_1289, opp(5) => n_1290, opp(4) => n_1291, 
                           opp(3) => n_1292, opp(2) => n_1293, opp(1) => n_1294
                           , opp(0) => n_1295);
   rast_addr_12_port <= '0';
   rast_addr_13_port <= '0';
   rast_addr_14_port <= '0';
   rast_addr_15_port <= '0';
   err <= '0';
   row_sel_1_port <= '0';

end SYN_struct;
