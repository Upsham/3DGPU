
module matrix_math_DW01_add_25 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] ,
         \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58;
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INVX1 U2 ( .A(n4), .Y(n5) );
  INVX1 U3 ( .A(n58), .Y(n6) );
  INVX1 U4 ( .A(n48), .Y(n1) );
  INVX2 U5 ( .A(n45), .Y(n48) );
  INVX2 U6 ( .A(n11), .Y(n34) );
  OR2X2 U7 ( .A(A[18]), .B(B[18]), .Y(n33) );
  XNOR2X1 U8 ( .A(n28), .B(n2), .Y(SUM[20]) );
  NAND2X1 U9 ( .A(n17), .B(n22), .Y(n2) );
  AND2X2 U10 ( .A(n52), .B(n58), .Y(SUM[14]) );
  INVX1 U11 ( .A(n4), .Y(n3) );
  INVX2 U12 ( .A(B[14]), .Y(n4) );
  OR2X1 U13 ( .A(n10), .B(n3), .Y(n52) );
  NAND2X1 U14 ( .A(n58), .B(n7), .Y(n8) );
  NAND2X1 U15 ( .A(n57), .B(n6), .Y(n9) );
  NAND2X1 U16 ( .A(n9), .B(n8), .Y(SUM[15]) );
  INVX1 U17 ( .A(n57), .Y(n7) );
  BUFX2 U18 ( .A(A[14]), .Y(n10) );
  AND2X2 U19 ( .A(n43), .B(n1), .Y(n11) );
  AND2X2 U20 ( .A(n11), .B(n33), .Y(n12) );
  XNOR2X1 U21 ( .A(n46), .B(n47), .Y(SUM[17]) );
  XNOR2X1 U22 ( .A(n38), .B(n39), .Y(SUM[18]) );
  XNOR2X1 U23 ( .A(n30), .B(n31), .Y(SUM[19]) );
  NAND2X1 U24 ( .A(n49), .B(n50), .Y(n25) );
  NAND2X1 U25 ( .A(n56), .B(n50), .Y(n54) );
  XOR2X1 U26 ( .A(n14), .B(n15), .Y(SUM[21]) );
  XOR2X1 U27 ( .A(B[21]), .B(A[21]), .Y(n15) );
  NAND2X1 U28 ( .A(n16), .B(n17), .Y(n14) );
  OAI21X1 U29 ( .A(n18), .B(n19), .C(n20), .Y(n16) );
  AND2X2 U30 ( .A(n21), .B(n22), .Y(n20) );
  NAND2X1 U31 ( .A(n23), .B(n24), .Y(n19) );
  NAND2X1 U32 ( .A(n12), .B(n25), .Y(n24) );
  NAND2X1 U33 ( .A(n26), .B(n27), .Y(n18) );
  OR2X2 U34 ( .A(A[20]), .B(B[20]), .Y(n22) );
  NAND2X1 U35 ( .A(B[20]), .B(A[20]), .Y(n17) );
  NAND2X1 U36 ( .A(n29), .B(n27), .Y(n28) );
  NAND2X1 U37 ( .A(n21), .B(n30), .Y(n29) );
  NAND2X1 U38 ( .A(n27), .B(n21), .Y(n31) );
  OR2X2 U39 ( .A(A[19]), .B(B[19]), .Y(n21) );
  NAND2X1 U40 ( .A(B[19]), .B(A[19]), .Y(n27) );
  NAND3X1 U41 ( .A(n23), .B(n26), .C(n32), .Y(n30) );
  NAND2X1 U42 ( .A(n25), .B(n12), .Y(n32) );
  NAND2X1 U43 ( .A(n35), .B(n33), .Y(n23) );
  NAND2X1 U44 ( .A(n36), .B(n37), .Y(n35) );
  NAND2X1 U45 ( .A(n26), .B(n33), .Y(n39) );
  NAND2X1 U46 ( .A(A[18]), .B(B[18]), .Y(n26) );
  OAI21X1 U47 ( .A(n40), .B(n34), .C(n41), .Y(n38) );
  AND2X2 U48 ( .A(n36), .B(n37), .Y(n41) );
  NAND2X1 U49 ( .A(n43), .B(n42), .Y(n36) );
  INVX2 U50 ( .A(n44), .Y(n42) );
  NAND2X1 U51 ( .A(n43), .B(n37), .Y(n47) );
  OR2X2 U52 ( .A(A[17]), .B(B[17]), .Y(n43) );
  NAND2X1 U53 ( .A(A[17]), .B(B[17]), .Y(n37) );
  OAI21X1 U54 ( .A(n40), .B(n48), .C(n44), .Y(n46) );
  INVX2 U55 ( .A(n25), .Y(n40) );
  NAND2X1 U56 ( .A(n51), .B(n53), .Y(n49) );
  AND2X2 U57 ( .A(B[14]), .B(A[14]), .Y(n53) );
  XNOR2X1 U58 ( .A(n54), .B(n55), .Y(SUM[16]) );
  NAND2X1 U59 ( .A(n45), .B(n44), .Y(n55) );
  NAND2X1 U60 ( .A(A[16]), .B(B[16]), .Y(n44) );
  OR2X2 U61 ( .A(B[16]), .B(A[16]), .Y(n45) );
  NAND2X1 U62 ( .A(n51), .B(n53), .Y(n56) );
  NAND2X1 U63 ( .A(n51), .B(n50), .Y(n57) );
  NAND2X1 U64 ( .A(A[15]), .B(B[15]), .Y(n50) );
  OR2X2 U65 ( .A(A[15]), .B(B[15]), .Y(n51) );
  NAND2X1 U66 ( .A(n5), .B(n10), .Y(n58) );
endmodule


module matrix_math_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][7] ,
         \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] ,
         \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] , \ab[2][13] ,
         \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][15] , \ab[1][14] ,
         \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] ,
         \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][14] , \ab[0][13] ,
         \ab[0][12] , \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] ,
         \ab[0][6] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[15][15] , \CARRYB[15][14] , \CARRYB[15][13] ,
         \CARRYB[15][12] , \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] ,
         \CARRYB[15][8] , \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] ,
         \CARRYB[15][4] , \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] ,
         \CARRYB[15][0] , \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][4] , \CARRYB[13][2] ,
         \CARRYB[13][1] , \CARRYB[13][0] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] ,
         \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][14] ,
         \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] ,
         \CARRYB[2][9] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][1] , \SUMB[15][15] , \SUMB[15][14] ,
         \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] ,
         \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] ,
         \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] ,
         \SUMB[15][1] , \SUMB[15][0] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] ,
         \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] ,
         \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][14] , \SUMB[12][13] ,
         \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] ,
         \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] , \SUMB[10][13] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] ,
         \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][14] , \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] ,
         \SUMB[3][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         ZA, ZB, \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] ,
         \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] ,
         \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] ,
         \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] ,
         \A1[1] , \A1[0] , \A2[22] , \A2[21] , \A2[14] , n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign ZA = A[15];
  assign ZB = B[15];

  FAX1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .C(\SUMB[14][9] ), .YC(
        \CARRYB[15][8] ), .YS(\SUMB[15][8] ) );
  FAX1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .C(\SUMB[14][10] ), .YC(
        \CARRYB[15][9] ), .YS(\SUMB[15][9] ) );
  FAX1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .C(\SUMB[14][11] ), 
        .YC(\CARRYB[15][10] ), .YS(\SUMB[15][10] ) );
  FAX1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .C(\SUMB[14][12] ), 
        .YC(\CARRYB[15][11] ), .YS(\SUMB[15][11] ) );
  FAX1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .C(\SUMB[14][13] ), 
        .YC(\CARRYB[15][12] ), .YS(\SUMB[15][12] ) );
  FAX1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .C(\SUMB[14][14] ), 
        .YC(\CARRYB[15][13] ), .YS(\SUMB[15][13] ) );
  FAX1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .C(\ab[14][15] ), .YC(
        \CARRYB[15][14] ), .YS(\SUMB[15][14] ) );
  FAX1 S14_15 ( .A(n1052), .B(n1051), .C(\ab[15][15] ), .YC(\CARRYB[15][15] ), 
        .YS(\SUMB[15][15] ) );
  FAX1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .C(\SUMB[13][10] ), 
        .YC(\CARRYB[14][9] ), .YS(\SUMB[14][9] ) );
  FAX1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .C(\SUMB[13][11] ), 
        .YC(\CARRYB[14][10] ), .YS(\SUMB[14][10] ) );
  FAX1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .C(\SUMB[13][12] ), 
        .YC(\CARRYB[14][11] ), .YS(\SUMB[14][11] ) );
  FAX1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .C(\SUMB[13][13] ), 
        .YC(\CARRYB[14][12] ), .YS(\SUMB[14][12] ) );
  FAX1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .C(\SUMB[13][14] ), 
        .YC(\CARRYB[14][13] ), .YS(\SUMB[14][13] ) );
  FAX1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .C(\ab[13][15] ), 
        .YC(\CARRYB[14][14] ), .YS(\SUMB[14][14] ) );
  FAX1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .C(\SUMB[12][10] ), 
        .YC(\CARRYB[13][9] ), .YS(\SUMB[13][9] ) );
  FAX1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .C(\SUMB[12][11] ), 
        .YC(\CARRYB[13][10] ), .YS(\SUMB[13][10] ) );
  FAX1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .C(\SUMB[12][12] ), 
        .YC(\CARRYB[13][11] ), .YS(\SUMB[13][11] ) );
  FAX1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .C(\SUMB[12][13] ), 
        .YC(\CARRYB[13][12] ), .YS(\SUMB[13][12] ) );
  FAX1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .C(\SUMB[12][14] ), 
        .YC(\CARRYB[13][13] ), .YS(\SUMB[13][13] ) );
  FAX1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .C(\ab[12][15] ), 
        .YC(\CARRYB[13][14] ), .YS(\SUMB[13][14] ) );
  FAX1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .C(\SUMB[11][12] ), 
        .YC(\CARRYB[12][11] ), .YS(\SUMB[12][11] ) );
  FAX1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .C(\SUMB[11][13] ), 
        .YC(\CARRYB[12][12] ), .YS(\SUMB[12][12] ) );
  FAX1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .C(\SUMB[11][14] ), 
        .YC(\CARRYB[12][13] ), .YS(\SUMB[12][13] ) );
  FAX1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .C(\ab[11][15] ), 
        .YC(\CARRYB[12][14] ), .YS(\SUMB[12][14] ) );
  FAX1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .C(\SUMB[10][2] ), .YC(
        \CARRYB[11][1] ), .YS(\SUMB[11][1] ) );
  FAX1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .C(\SUMB[10][10] ), 
        .YC(\CARRYB[11][9] ), .YS(\SUMB[11][9] ) );
  FAX1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .C(\SUMB[10][13] ), 
        .YC(\CARRYB[11][12] ), .YS(\SUMB[11][12] ) );
  FAX1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .C(\SUMB[10][14] ), 
        .YC(\CARRYB[11][13] ), .YS(\SUMB[11][13] ) );
  FAX1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .C(\ab[10][15] ), 
        .YC(\CARRYB[11][14] ), .YS(\SUMB[11][14] ) );
  FAX1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .C(\SUMB[9][13] ), 
        .YC(\CARRYB[10][12] ), .YS(\SUMB[10][12] ) );
  FAX1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .C(\SUMB[9][14] ), 
        .YC(\CARRYB[10][13] ), .YS(\SUMB[10][13] ) );
  FAX1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .C(\ab[9][15] ), .YC(
        \CARRYB[10][14] ), .YS(\SUMB[10][14] ) );
  FAX1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .C(\SUMB[8][1] ), .YC(
        \CARRYB[9][0] ), .YS(\A1[7] ) );
  FAX1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .C(\SUMB[8][14] ), .YC(
        \CARRYB[9][13] ), .YS(\SUMB[9][13] ) );
  FAX1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .C(\ab[8][15] ), .YC(
        \CARRYB[9][14] ), .YS(\SUMB[9][14] ) );
  FAX1 S2_8_13 ( .A(\ab[8][13] ), .B(\SUMB[7][14] ), .C(\CARRYB[7][13] ), .YC(
        \CARRYB[8][13] ), .YS(\SUMB[8][13] ) );
  FAX1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .C(\ab[7][15] ), .YC(
        \CARRYB[8][14] ), .YS(\SUMB[8][14] ) );
  FAX1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .C(\ab[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_6_12 ( .A(\ab[6][12] ), .B(n286), .C(\SUMB[5][13] ), .YC(
        \CARRYB[6][12] ), .YS(\SUMB[6][12] ) );
  FAX1 S2_6_13 ( .A(\ab[6][13] ), .B(n242), .C(\SUMB[5][14] ), .YC(
        \CARRYB[6][13] ), .YS(\SUMB[6][13] ) );
  FAX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .C(\SUMB[4][13] ), .YC(
        \CARRYB[5][12] ), .YS(\SUMB[5][12] ) );
  FAX1 S2_5_13 ( .A(\ab[5][13] ), .B(n367), .C(\SUMB[4][14] ), .YC(
        \CARRYB[5][13] ), .YS(\SUMB[5][13] ) );
  FAX1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .C(\ab[4][15] ), .YC(
        \CARRYB[5][14] ), .YS(\SUMB[5][14] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .C(\SUMB[3][14] ), .YC(
        \CARRYB[4][13] ), .YS(\SUMB[4][13] ) );
  FAX1 S1_3_0 ( .A(\ab[3][0] ), .B(n968), .C(\SUMB[2][1] ), .YC(\CARRYB[3][0] ), .YS(\A1[1] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n958), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .C(\SUMB[1][2] ), .YC(
        \CARRYB[2][1] ), .YS(\SUMB[2][1] ) );
  matrix_math_DW01_add_25 FS_1 ( .A({n1050, \A1[28] , \A1[27] , \A1[26] , 
        \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , 
        \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n72, n71, n70, n69, 
        n68, n67, n66, \A2[22] , \A2[21] , n957, n956, n954, n952, n953, n955, 
        \A2[14] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, PRODUCT[23:2]}) );
  XOR2X1 U2 ( .A(n3), .B(\ab[0][10] ), .Y(\SUMB[1][9] ) );
  AND2X2 U3 ( .A(n423), .B(B[9]), .Y(n3) );
  INVX2 U4 ( .A(n1019), .Y(n4) );
  INVX2 U5 ( .A(n1019), .Y(n5) );
  INVX2 U6 ( .A(n1019), .Y(n1020) );
  INVX2 U7 ( .A(A[2]), .Y(n1019) );
  INVX4 U8 ( .A(n1017), .Y(n423) );
  INVX1 U9 ( .A(\SUMB[2][7] ), .Y(n323) );
  XNOR2X1 U10 ( .A(n282), .B(n41), .Y(n6) );
  INVX2 U11 ( .A(n8), .Y(n9) );
  NAND3X1 U12 ( .A(n259), .B(n258), .C(n260), .Y(n7) );
  INVX1 U13 ( .A(n1018), .Y(n8) );
  BUFX2 U14 ( .A(n5), .Y(n10) );
  NAND3X1 U15 ( .A(n335), .B(n336), .C(n337), .Y(n11) );
  BUFX2 U16 ( .A(n418), .Y(n12) );
  XOR2X1 U17 ( .A(\CARRYB[6][6] ), .B(n13), .Y(n19) );
  INVX8 U18 ( .A(\ab[7][6] ), .Y(n13) );
  NAND3X1 U19 ( .A(n511), .B(n510), .C(n509), .Y(n14) );
  NAND3X1 U20 ( .A(n455), .B(n454), .C(n456), .Y(n15) );
  XOR2X1 U21 ( .A(n16), .B(n373), .Y(\SUMB[8][4] ) );
  INVX1 U22 ( .A(\SUMB[7][5] ), .Y(n16) );
  XNOR2X1 U23 ( .A(n17), .B(\SUMB[4][7] ), .Y(\SUMB[5][6] ) );
  XNOR2X1 U24 ( .A(\CARRYB[4][6] ), .B(\ab[5][6] ), .Y(n17) );
  BUFX2 U25 ( .A(\SUMB[5][11] ), .Y(n18) );
  INVX2 U26 ( .A(A[0]), .Y(n1016) );
  XOR2X1 U27 ( .A(n374), .B(n19), .Y(\SUMB[7][6] ) );
  NAND3X1 U28 ( .A(n746), .B(n747), .C(n748), .Y(n20) );
  AND2X1 U29 ( .A(n423), .B(B[9]), .Y(\ab[1][9] ) );
  INVX1 U30 ( .A(\SUMB[14][6] ), .Y(n21) );
  INVX1 U31 ( .A(n21), .Y(n22) );
  XOR2X1 U32 ( .A(\CARRYB[13][2] ), .B(n23), .Y(n315) );
  INVX8 U33 ( .A(\ab[14][2] ), .Y(n23) );
  XNOR2X1 U34 ( .A(n24), .B(n174), .Y(\SUMB[4][5] ) );
  XOR2X1 U35 ( .A(n407), .B(\ab[4][5] ), .Y(n24) );
  XNOR2X1 U36 ( .A(\CARRYB[14][0] ), .B(n25), .Y(n302) );
  INVX8 U37 ( .A(\ab[15][0] ), .Y(n25) );
  BUFX4 U38 ( .A(\ab[2][12] ), .Y(n160) );
  XOR2X1 U39 ( .A(\SUMB[15][3] ), .B(\CARRYB[15][2] ), .Y(\A1[16] ) );
  INVX1 U40 ( .A(\CARRYB[15][2] ), .Y(n593) );
  XNOR2X1 U41 ( .A(n26), .B(n347), .Y(\SUMB[10][2] ) );
  XOR2X1 U42 ( .A(\CARRYB[9][2] ), .B(\ab[10][2] ), .Y(n26) );
  XOR2X1 U43 ( .A(n134), .B(n27), .Y(n504) );
  INVX8 U44 ( .A(\ab[14][3] ), .Y(n27) );
  XOR2X1 U45 ( .A(n229), .B(n29), .Y(n28) );
  XOR2X1 U46 ( .A(n229), .B(n29), .Y(\SUMB[12][3] ) );
  AND2X2 U47 ( .A(n766), .B(n102), .Y(n29) );
  AND2X2 U48 ( .A(n984), .B(\ab[1][14] ), .Y(n30) );
  XNOR2X1 U49 ( .A(n31), .B(\CARRYB[11][8] ), .Y(n642) );
  INVX8 U50 ( .A(\ab[12][8] ), .Y(n31) );
  AND2X1 U51 ( .A(\SUMB[15][6] ), .B(\CARRYB[15][5] ), .Y(n957) );
  XNOR2X1 U52 ( .A(n32), .B(n33), .Y(\SUMB[9][5] ) );
  XNOR2X1 U53 ( .A(\CARRYB[8][5] ), .B(\ab[9][5] ), .Y(n32) );
  XOR2X1 U54 ( .A(n447), .B(n448), .Y(n33) );
  XOR2X1 U55 ( .A(n34), .B(\SUMB[10][7] ), .Y(\SUMB[11][6] ) );
  XOR2X1 U56 ( .A(\CARRYB[10][6] ), .B(\ab[11][6] ), .Y(n34) );
  XNOR2X1 U57 ( .A(n508), .B(n35), .Y(\SUMB[6][4] ) );
  INVX1 U58 ( .A(\SUMB[5][5] ), .Y(n35) );
  XNOR2X1 U59 ( .A(\SUMB[8][4] ), .B(n36), .Y(\SUMB[9][3] ) );
  XNOR2X1 U60 ( .A(\CARRYB[8][3] ), .B(\ab[9][3] ), .Y(n36) );
  XOR2X1 U61 ( .A(n37), .B(n415), .Y(\SUMB[2][8] ) );
  XOR2X1 U62 ( .A(\SUMB[1][9] ), .B(\ab[2][8] ), .Y(n37) );
  XOR2X1 U63 ( .A(n38), .B(\ab[10][1] ), .Y(n40) );
  INVX1 U64 ( .A(\SUMB[9][2] ), .Y(n38) );
  XOR2X1 U65 ( .A(n39), .B(n40), .Y(\SUMB[10][1] ) );
  INVX1 U66 ( .A(n7), .Y(n39) );
  XOR2X1 U67 ( .A(\SUMB[6][10] ), .B(n107), .Y(n41) );
  XNOR2X1 U68 ( .A(n42), .B(\SUMB[3][11] ), .Y(\SUMB[4][10] ) );
  XNOR2X1 U69 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .Y(n42) );
  XOR2X1 U70 ( .A(n43), .B(\SUMB[8][9] ), .Y(\SUMB[9][8] ) );
  XNOR2X1 U71 ( .A(n248), .B(\CARRYB[8][8] ), .Y(n43) );
  NAND3X1 U72 ( .A(n483), .B(n482), .C(n484), .Y(n44) );
  NAND3X1 U73 ( .A(n865), .B(n866), .C(n867), .Y(n45) );
  INVX1 U74 ( .A(\SUMB[15][4] ), .Y(n46) );
  INVX1 U75 ( .A(n46), .Y(n47) );
  BUFX4 U76 ( .A(n1016), .Y(n655) );
  NAND3X1 U77 ( .A(n561), .B(n560), .C(n562), .Y(n48) );
  NAND3X1 U78 ( .A(n156), .B(n155), .C(n157), .Y(n49) );
  NAND3X1 U79 ( .A(n939), .B(n940), .C(n941), .Y(n50) );
  NAND3X1 U80 ( .A(n546), .B(n545), .C(n547), .Y(n51) );
  BUFX2 U81 ( .A(\CARRYB[9][0] ), .Y(n52) );
  BUFX2 U82 ( .A(\CARRYB[6][1] ), .Y(n53) );
  NAND3X1 U83 ( .A(n856), .B(n857), .C(n858), .Y(n54) );
  NAND3X1 U84 ( .A(n805), .B(n806), .C(n807), .Y(n55) );
  NAND3X1 U85 ( .A(n574), .B(n572), .C(n573), .Y(n56) );
  NAND3X1 U86 ( .A(n379), .B(n378), .C(n380), .Y(n57) );
  XNOR2X1 U87 ( .A(\CARRYB[7][6] ), .B(n58), .Y(n447) );
  INVX8 U88 ( .A(n104), .Y(n58) );
  INVX4 U89 ( .A(n989), .Y(n974) );
  INVX4 U90 ( .A(B[0]), .Y(n989) );
  AND2X2 U91 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n59) );
  NAND3X1 U92 ( .A(n492), .B(n493), .C(n494), .Y(n60) );
  XOR2X1 U93 ( .A(n61), .B(n62), .Y(\SUMB[11][4] ) );
  XNOR2X1 U94 ( .A(n970), .B(\ab[11][4] ), .Y(n61) );
  XNOR2X1 U95 ( .A(n220), .B(n444), .Y(n62) );
  INVX2 U96 ( .A(\SUMB[12][2] ), .Y(n400) );
  INVX2 U97 ( .A(\SUMB[2][6] ), .Y(n385) );
  XOR2X1 U98 ( .A(\CARRYB[14][3] ), .B(n63), .Y(n595) );
  INVX8 U99 ( .A(\ab[15][3] ), .Y(n63) );
  XNOR2X1 U100 ( .A(n64), .B(\SUMB[10][6] ), .Y(\SUMB[11][5] ) );
  XNOR2X1 U101 ( .A(\CARRYB[10][5] ), .B(\ab[11][5] ), .Y(n64) );
  INVX2 U102 ( .A(\SUMB[6][7] ), .Y(n374) );
  INVX2 U103 ( .A(\SUMB[12][4] ), .Y(n221) );
  XNOR2X1 U104 ( .A(n65), .B(\SUMB[3][10] ), .Y(\SUMB[4][9] ) );
  XNOR2X1 U105 ( .A(n325), .B(\ab[4][9] ), .Y(n65) );
  INVX1 U106 ( .A(n970), .Y(n971) );
  INVX2 U107 ( .A(\ab[8][8] ), .Y(n280) );
  INVX2 U108 ( .A(\ab[9][7] ), .Y(n200) );
  INVX2 U109 ( .A(n414), .Y(n178) );
  INVX2 U110 ( .A(\ab[5][9] ), .Y(n530) );
  INVX2 U111 ( .A(\ab[3][12] ), .Y(n150) );
  INVX2 U112 ( .A(\ab[6][9] ), .Y(n149) );
  INVX2 U113 ( .A(\ab[10][5] ), .Y(n130) );
  INVX2 U114 ( .A(\ab[9][8] ), .Y(n248) );
  INVX2 U115 ( .A(B[4]), .Y(n997) );
  INVX2 U116 ( .A(\ab[13][5] ), .Y(n201) );
  INVX2 U117 ( .A(\ab[12][7] ), .Y(n568) );
  INVX2 U118 ( .A(\ab[5][8] ), .Y(n362) );
  INVX2 U119 ( .A(\ab[6][8] ), .Y(n162) );
  INVX2 U120 ( .A(\ab[4][6] ), .Y(n317) );
  INVX2 U121 ( .A(\ab[3][5] ), .Y(n250) );
  INVX2 U122 ( .A(\ab[2][15] ), .Y(n243) );
  INVX2 U123 ( .A(\ab[8][6] ), .Y(n104) );
  INVX2 U124 ( .A(\ab[5][10] ), .Y(n279) );
  INVX2 U125 ( .A(\ab[4][3] ), .Y(n501) );
  INVX2 U126 ( .A(\ab[8][4] ), .Y(n175) );
  INVX2 U127 ( .A(\ab[12][3] ), .Y(n222) );
  INVX2 U128 ( .A(\ab[6][10] ), .Y(n247) );
  INVX2 U129 ( .A(\ab[15][2] ), .Y(n476) );
  INVX1 U130 ( .A(\SUMB[6][14] ), .Y(n296) );
  INVX2 U131 ( .A(\ab[15][4] ), .Y(n210) );
  INVX2 U132 ( .A(\ab[12][1] ), .Y(n804) );
  INVX2 U133 ( .A(\CARRYB[15][6] ), .Y(n294) );
  INVX2 U134 ( .A(B[11]), .Y(n1008) );
  INVX4 U135 ( .A(n1010), .Y(n1011) );
  INVX2 U136 ( .A(B[14]), .Y(n1014) );
  AND2X2 U137 ( .A(\SUMB[15][9] ), .B(\CARRYB[15][8] ), .Y(n66) );
  AND2X2 U138 ( .A(\SUMB[15][10] ), .B(\CARRYB[15][9] ), .Y(n67) );
  AND2X2 U139 ( .A(\SUMB[15][11] ), .B(\CARRYB[15][10] ), .Y(n68) );
  AND2X2 U140 ( .A(\SUMB[15][12] ), .B(\CARRYB[15][11] ), .Y(n69) );
  AND2X2 U141 ( .A(\SUMB[15][13] ), .B(\CARRYB[15][12] ), .Y(n70) );
  AND2X2 U142 ( .A(\SUMB[15][14] ), .B(\CARRYB[15][13] ), .Y(n71) );
  AND2X2 U143 ( .A(\SUMB[15][15] ), .B(\CARRYB[15][14] ), .Y(n72) );
  INVX1 U144 ( .A(\CARRYB[3][1] ), .Y(n988) );
  INVX1 U145 ( .A(\CARRYB[6][13] ), .Y(n368) );
  AND2X2 U146 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(n73) );
  INVX2 U147 ( .A(n959), .Y(n979) );
  INVX2 U148 ( .A(B[10]), .Y(n1006) );
  INVX2 U149 ( .A(\ab[13][3] ), .Y(n477) );
  XOR2X1 U150 ( .A(n412), .B(n74), .Y(\SUMB[8][1] ) );
  XNOR2X1 U151 ( .A(\CARRYB[7][1] ), .B(\ab[8][1] ), .Y(n74) );
  BUFX2 U152 ( .A(\SUMB[4][4] ), .Y(n75) );
  BUFX2 U153 ( .A(\SUMB[13][2] ), .Y(n76) );
  BUFX2 U154 ( .A(\SUMB[4][11] ), .Y(n77) );
  BUFX2 U155 ( .A(\CARRYB[3][2] ), .Y(n78) );
  XOR2X1 U156 ( .A(n143), .B(n92), .Y(n79) );
  XNOR2X1 U157 ( .A(n80), .B(\ab[0][14] ), .Y(\SUMB[1][13] ) );
  NAND2X1 U158 ( .A(n1018), .B(n1013), .Y(n80) );
  BUFX2 U159 ( .A(\SUMB[8][2] ), .Y(n81) );
  NAND3X1 U160 ( .A(n709), .B(n710), .C(n711), .Y(n82) );
  XNOR2X1 U161 ( .A(n83), .B(\SUMB[12][6] ), .Y(\SUMB[13][5] ) );
  XOR2X1 U162 ( .A(\CARRYB[12][5] ), .B(n201), .Y(n83) );
  XNOR2X1 U163 ( .A(n84), .B(\CARRYB[5][9] ), .Y(\SUMB[6][9] ) );
  XOR2X1 U164 ( .A(\SUMB[5][10] ), .B(n149), .Y(n84) );
  BUFX2 U165 ( .A(\CARRYB[7][0] ), .Y(n85) );
  BUFX2 U166 ( .A(\SUMB[7][1] ), .Y(n86) );
  NAND3X1 U167 ( .A(n839), .B(n838), .C(n840), .Y(n87) );
  NAND3X1 U168 ( .A(n781), .B(n782), .C(n783), .Y(n88) );
  XOR2X1 U169 ( .A(n315), .B(n442), .Y(n89) );
  INVX2 U170 ( .A(\SUMB[13][3] ), .Y(n442) );
  XOR2X1 U171 ( .A(n90), .B(\SUMB[6][9] ), .Y(\SUMB[7][8] ) );
  XOR2X1 U172 ( .A(\CARRYB[6][8] ), .B(\ab[7][8] ), .Y(n90) );
  XNOR2X1 U173 ( .A(\CARRYB[8][6] ), .B(\ab[9][6] ), .Y(n148) );
  BUFX2 U174 ( .A(n864), .Y(n91) );
  BUFX2 U175 ( .A(\CARRYB[9][4] ), .Y(n92) );
  NAND3X1 U176 ( .A(n868), .B(n869), .C(n870), .Y(n93) );
  NAND3X1 U177 ( .A(n541), .B(n542), .C(n540), .Y(n94) );
  NAND3X1 U178 ( .A(n659), .B(n660), .C(n661), .Y(n95) );
  NOR2X1 U179 ( .A(n1012), .B(n655), .Y(n96) );
  NAND3X1 U180 ( .A(n827), .B(n828), .C(n829), .Y(n97) );
  BUFX2 U181 ( .A(\SUMB[2][5] ), .Y(n98) );
  XNOR2X1 U182 ( .A(n99), .B(n59), .Y(\SUMB[2][5] ) );
  XNOR2X1 U183 ( .A(\SUMB[1][6] ), .B(\ab[2][5] ), .Y(n99) );
  XOR2X1 U184 ( .A(n100), .B(n385), .Y(\SUMB[3][5] ) );
  XOR2X1 U185 ( .A(\CARRYB[2][5] ), .B(n250), .Y(n100) );
  NAND2X1 U186 ( .A(n765), .B(n767), .Y(n101) );
  INVX2 U187 ( .A(n101), .Y(n102) );
  INVX2 U188 ( .A(\CARRYB[15][4] ), .Y(n293) );
  XOR2X1 U189 ( .A(n103), .B(n158), .Y(\SUMB[5][5] ) );
  XNOR2X1 U190 ( .A(\CARRYB[4][5] ), .B(\ab[5][5] ), .Y(n103) );
  XNOR2X1 U191 ( .A(n105), .B(\SUMB[11][5] ), .Y(\SUMB[12][4] ) );
  XNOR2X1 U192 ( .A(\CARRYB[11][4] ), .B(\ab[12][4] ), .Y(n105) );
  BUFX2 U193 ( .A(\SUMB[3][9] ), .Y(n106) );
  XOR2X1 U194 ( .A(\CARRYB[6][9] ), .B(\ab[7][9] ), .Y(n107) );
  XOR2X1 U195 ( .A(\SUMB[6][10] ), .B(n107), .Y(\SUMB[7][9] ) );
  NAND2X1 U196 ( .A(\SUMB[6][10] ), .B(\CARRYB[6][9] ), .Y(n108) );
  NAND2X1 U197 ( .A(\SUMB[6][10] ), .B(\ab[7][9] ), .Y(n109) );
  NAND2X1 U198 ( .A(\CARRYB[6][9] ), .B(\ab[7][9] ), .Y(n110) );
  NAND3X1 U199 ( .A(n109), .B(n108), .C(n110), .Y(\CARRYB[7][9] ) );
  NAND3X1 U200 ( .A(n821), .B(n822), .C(n823), .Y(n111) );
  NAND3X1 U201 ( .A(n818), .B(n819), .C(n820), .Y(n112) );
  XOR2X1 U202 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .Y(n113) );
  XOR2X1 U203 ( .A(n113), .B(\SUMB[13][9] ), .Y(\SUMB[14][8] ) );
  XOR2X1 U204 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .Y(n114) );
  XOR2X1 U205 ( .A(n114), .B(\SUMB[14][8] ), .Y(\SUMB[15][7] ) );
  NAND2X1 U206 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .Y(n115) );
  NAND2X1 U207 ( .A(\ab[14][8] ), .B(\SUMB[13][9] ), .Y(n116) );
  NAND2X1 U208 ( .A(\CARRYB[13][8] ), .B(\SUMB[13][9] ), .Y(n117) );
  NAND3X1 U209 ( .A(n115), .B(n116), .C(n117), .Y(\CARRYB[14][8] ) );
  NAND2X1 U210 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .Y(n118) );
  NAND2X1 U211 ( .A(\ab[15][7] ), .B(\SUMB[14][8] ), .Y(n119) );
  NAND2X1 U212 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Y(n120) );
  NAND3X1 U213 ( .A(n118), .B(n119), .C(n120), .Y(\CARRYB[15][7] ) );
  XOR2X1 U214 ( .A(\SUMB[8][11] ), .B(\ab[9][10] ), .Y(n121) );
  XOR2X1 U215 ( .A(n121), .B(\CARRYB[8][10] ), .Y(\SUMB[9][10] ) );
  NAND2X1 U216 ( .A(\CARRYB[8][10] ), .B(\SUMB[8][11] ), .Y(n122) );
  NAND2X1 U217 ( .A(\CARRYB[8][10] ), .B(\ab[9][10] ), .Y(n123) );
  NAND2X1 U218 ( .A(\SUMB[8][11] ), .B(\ab[9][10] ), .Y(n124) );
  NAND3X1 U219 ( .A(n123), .B(n122), .C(n124), .Y(\CARRYB[9][10] ) );
  XOR2X1 U220 ( .A(\CARRYB[12][8] ), .B(\ab[13][8] ), .Y(n125) );
  XOR2X1 U221 ( .A(\SUMB[12][9] ), .B(n125), .Y(\SUMB[13][8] ) );
  NAND2X1 U222 ( .A(\SUMB[12][9] ), .B(\CARRYB[12][8] ), .Y(n126) );
  NAND2X1 U223 ( .A(\SUMB[12][9] ), .B(\ab[13][8] ), .Y(n127) );
  NAND2X1 U224 ( .A(\CARRYB[12][8] ), .B(\ab[13][8] ), .Y(n128) );
  NAND3X1 U225 ( .A(n127), .B(n126), .C(n128), .Y(\CARRYB[13][8] ) );
  NAND3X1 U226 ( .A(n916), .B(n915), .C(n917), .Y(n129) );
  XNOR2X1 U227 ( .A(\CARRYB[9][5] ), .B(n130), .Y(n220) );
  XOR2X1 U228 ( .A(n131), .B(n179), .Y(\SUMB[6][2] ) );
  XOR2X1 U229 ( .A(\ab[6][2] ), .B(n50), .Y(n131) );
  INVX4 U230 ( .A(n991), .Y(n980) );
  INVX2 U231 ( .A(n1016), .Y(n401) );
  INVX1 U232 ( .A(n593), .Y(n132) );
  XNOR2X1 U233 ( .A(n504), .B(n254), .Y(n133) );
  NAND3X1 U234 ( .A(n845), .B(n847), .C(n846), .Y(n134) );
  XNOR2X1 U235 ( .A(n135), .B(n136), .Y(\SUMB[12][2] ) );
  XOR2X1 U236 ( .A(\CARRYB[11][2] ), .B(\ab[12][2] ), .Y(n135) );
  INVX1 U237 ( .A(\SUMB[11][3] ), .Y(n136) );
  BUFX2 U238 ( .A(\SUMB[8][3] ), .Y(n137) );
  XNOR2X1 U239 ( .A(n138), .B(\SUMB[7][4] ), .Y(\SUMB[8][3] ) );
  XNOR2X1 U240 ( .A(\CARRYB[7][3] ), .B(\ab[8][3] ), .Y(n138) );
  AND2X2 U241 ( .A(n1018), .B(n1013), .Y(n139) );
  XOR2X1 U242 ( .A(n140), .B(n221), .Y(\SUMB[13][3] ) );
  XOR2X1 U243 ( .A(\CARRYB[12][3] ), .B(n477), .Y(n140) );
  XOR2X1 U244 ( .A(n141), .B(n142), .Y(\SUMB[7][3] ) );
  XNOR2X1 U245 ( .A(\CARRYB[6][3] ), .B(\ab[7][3] ), .Y(n141) );
  INVX1 U246 ( .A(\SUMB[6][4] ), .Y(n142) );
  XOR2X1 U247 ( .A(\SUMB[9][5] ), .B(\ab[10][4] ), .Y(n143) );
  XOR2X1 U248 ( .A(n143), .B(n92), .Y(\SUMB[10][4] ) );
  NAND2X1 U249 ( .A(\SUMB[9][5] ), .B(\CARRYB[9][4] ), .Y(n144) );
  NAND2X1 U250 ( .A(\CARRYB[9][4] ), .B(\ab[10][4] ), .Y(n145) );
  NAND2X1 U251 ( .A(\SUMB[9][5] ), .B(\ab[10][4] ), .Y(n146) );
  NAND3X1 U252 ( .A(n145), .B(n146), .C(n144), .Y(\CARRYB[10][4] ) );
  XOR2X1 U253 ( .A(n148), .B(n147), .Y(\SUMB[9][6] ) );
  INVX2 U254 ( .A(\SUMB[8][7] ), .Y(n147) );
  INVX4 U255 ( .A(n1006), .Y(n1007) );
  XOR2X1 U256 ( .A(\CARRYB[2][12] ), .B(n150), .Y(n151) );
  XNOR2X1 U257 ( .A(n151), .B(\SUMB[2][13] ), .Y(\SUMB[3][12] ) );
  INVX2 U258 ( .A(\CARRYB[7][9] ), .Y(n289) );
  XNOR2X1 U259 ( .A(\ab[1][10] ), .B(n152), .Y(\SUMB[1][10] ) );
  NAND2X1 U260 ( .A(n1009), .B(n401), .Y(n152) );
  XOR2X1 U261 ( .A(\CARRYB[4][7] ), .B(\ab[5][7] ), .Y(n771) );
  XNOR2X1 U262 ( .A(n153), .B(n465), .Y(\SUMB[2][9] ) );
  XOR2X1 U263 ( .A(\ab[2][9] ), .B(n760), .Y(n153) );
  NAND3X1 U264 ( .A(n266), .B(n265), .C(n267), .Y(n154) );
  AND2X2 U265 ( .A(\CARRYB[15][3] ), .B(n47), .Y(n954) );
  NAND2X1 U266 ( .A(\SUMB[8][4] ), .B(n57), .Y(n155) );
  NAND2X1 U267 ( .A(\SUMB[8][4] ), .B(\ab[9][3] ), .Y(n156) );
  NAND2X1 U268 ( .A(n57), .B(\ab[9][3] ), .Y(n157) );
  NAND3X1 U269 ( .A(n156), .B(n155), .C(n157), .Y(\CARRYB[9][3] ) );
  INVX2 U270 ( .A(\SUMB[4][6] ), .Y(n158) );
  NAND3X1 U271 ( .A(n656), .B(n657), .C(n658), .Y(n159) );
  BUFX2 U272 ( .A(n903), .Y(n161) );
  XOR2X1 U273 ( .A(\CARRYB[7][7] ), .B(\ab[8][7] ), .Y(n575) );
  XOR2X1 U274 ( .A(\CARRYB[5][8] ), .B(n162), .Y(n307) );
  BUFX2 U275 ( .A(n1009), .Y(n163) );
  INVX4 U276 ( .A(n1008), .Y(n1009) );
  NAND3X1 U277 ( .A(n311), .B(n310), .C(n312), .Y(n164) );
  NAND3X1 U278 ( .A(n436), .B(n437), .C(n438), .Y(n165) );
  XNOR2X1 U279 ( .A(n166), .B(n167), .Y(\SUMB[6][6] ) );
  XOR2X1 U280 ( .A(\SUMB[5][7] ), .B(\ab[6][6] ), .Y(n166) );
  INVX1 U281 ( .A(\CARRYB[5][6] ), .Y(n167) );
  XNOR2X1 U282 ( .A(n883), .B(n168), .Y(\SUMB[12][1] ) );
  INVX2 U283 ( .A(\SUMB[11][2] ), .Y(n168) );
  XOR2X1 U284 ( .A(\CARRYB[6][10] ), .B(\ab[7][10] ), .Y(n169) );
  XOR2X1 U285 ( .A(\SUMB[6][11] ), .B(n169), .Y(\SUMB[7][10] ) );
  NAND2X1 U286 ( .A(\SUMB[6][11] ), .B(n54), .Y(n170) );
  NAND2X1 U287 ( .A(\SUMB[6][11] ), .B(\ab[7][10] ), .Y(n171) );
  NAND2X1 U288 ( .A(n54), .B(\ab[7][10] ), .Y(n172) );
  NAND3X1 U289 ( .A(n171), .B(n170), .C(n172), .Y(\CARRYB[7][10] ) );
  XNOR2X1 U290 ( .A(n173), .B(n240), .Y(\SUMB[4][6] ) );
  XNOR2X1 U291 ( .A(n841), .B(n317), .Y(n173) );
  INVX1 U292 ( .A(\SUMB[3][6] ), .Y(n174) );
  XOR2X1 U293 ( .A(\CARRYB[7][4] ), .B(n175), .Y(n373) );
  BUFX2 U294 ( .A(\SUMB[2][2] ), .Y(n176) );
  INVX2 U295 ( .A(n182), .Y(n183) );
  XNOR2X1 U296 ( .A(n177), .B(\SUMB[13][7] ), .Y(\SUMB[14][6] ) );
  XNOR2X1 U297 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .Y(n177) );
  XOR2X1 U298 ( .A(n460), .B(n178), .Y(n219) );
  BUFX2 U299 ( .A(\SUMB[5][3] ), .Y(n179) );
  NAND3X1 U300 ( .A(n936), .B(n937), .C(n938), .Y(n180) );
  INVX2 U301 ( .A(\ab[2][7] ), .Y(n381) );
  AND2X2 U302 ( .A(n1009), .B(n402), .Y(n181) );
  INVX1 U303 ( .A(n802), .Y(n182) );
  XOR2X1 U304 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .Y(n184) );
  XOR2X1 U305 ( .A(n184), .B(\SUMB[10][12] ), .Y(\SUMB[11][11] ) );
  XOR2X1 U306 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .Y(n185) );
  XOR2X1 U307 ( .A(n185), .B(\SUMB[11][11] ), .Y(\SUMB[12][10] ) );
  NAND2X1 U308 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .Y(n186) );
  NAND2X1 U309 ( .A(\ab[11][11] ), .B(\SUMB[10][12] ), .Y(n187) );
  NAND2X1 U310 ( .A(\CARRYB[10][11] ), .B(\SUMB[10][12] ), .Y(n188) );
  NAND3X1 U311 ( .A(n186), .B(n187), .C(n188), .Y(\CARRYB[11][11] ) );
  NAND2X1 U312 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .Y(n189) );
  NAND2X1 U313 ( .A(\ab[12][10] ), .B(\SUMB[11][11] ), .Y(n190) );
  NAND2X1 U314 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Y(n191) );
  NAND3X1 U315 ( .A(n189), .B(n190), .C(n191), .Y(\CARRYB[12][10] ) );
  XOR2X1 U316 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .Y(n192) );
  XOR2X1 U317 ( .A(n192), .B(\SUMB[8][13] ), .Y(\SUMB[9][12] ) );
  XOR2X1 U318 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .Y(n193) );
  XOR2X1 U319 ( .A(n193), .B(\SUMB[9][12] ), .Y(\SUMB[10][11] ) );
  NAND2X1 U320 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .Y(n194) );
  NAND2X1 U321 ( .A(\ab[9][12] ), .B(\SUMB[8][13] ), .Y(n195) );
  NAND2X1 U322 ( .A(\CARRYB[8][12] ), .B(\SUMB[8][13] ), .Y(n196) );
  NAND3X1 U323 ( .A(n194), .B(n195), .C(n196), .Y(\CARRYB[9][12] ) );
  NAND2X1 U324 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .Y(n197) );
  NAND2X1 U325 ( .A(\ab[10][11] ), .B(\SUMB[9][12] ), .Y(n198) );
  NAND2X1 U326 ( .A(\CARRYB[9][11] ), .B(\SUMB[9][12] ), .Y(n199) );
  NAND3X1 U327 ( .A(n197), .B(n198), .C(n199), .Y(\CARRYB[10][11] ) );
  XOR2X1 U328 ( .A(\CARRYB[3][11] ), .B(\ab[4][11] ), .Y(n281) );
  XOR2X1 U329 ( .A(\CARRYB[8][7] ), .B(n200), .Y(n274) );
  XOR2X1 U330 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .Y(n202) );
  XOR2X1 U331 ( .A(n202), .B(\SUMB[10][11] ), .Y(\SUMB[11][10] ) );
  XOR2X1 U332 ( .A(\ab[12][9] ), .B(n216), .Y(n203) );
  XOR2X1 U333 ( .A(n203), .B(\SUMB[11][10] ), .Y(\SUMB[12][9] ) );
  NAND2X1 U334 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .Y(n204) );
  NAND2X1 U335 ( .A(\ab[11][10] ), .B(\SUMB[10][11] ), .Y(n205) );
  NAND2X1 U336 ( .A(\CARRYB[10][10] ), .B(\SUMB[10][11] ), .Y(n206) );
  NAND3X1 U337 ( .A(n204), .B(n205), .C(n206), .Y(\CARRYB[11][10] ) );
  NAND2X1 U338 ( .A(\ab[12][9] ), .B(n216), .Y(n207) );
  NAND2X1 U339 ( .A(\ab[12][9] ), .B(\SUMB[11][10] ), .Y(n208) );
  NAND2X1 U340 ( .A(n216), .B(\SUMB[11][10] ), .Y(n209) );
  NAND3X1 U341 ( .A(n207), .B(n208), .C(n209), .Y(\CARRYB[12][9] ) );
  XNOR2X1 U342 ( .A(\CARRYB[14][4] ), .B(n210), .Y(n741) );
  XOR2X1 U343 ( .A(n211), .B(n212), .Y(\SUMB[7][11] ) );
  XNOR2X1 U344 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .Y(n211) );
  INVX1 U345 ( .A(\SUMB[6][12] ), .Y(n212) );
  XNOR2X1 U346 ( .A(n213), .B(\SUMB[8][12] ), .Y(\SUMB[9][11] ) );
  XNOR2X1 U347 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .Y(n213) );
  NAND3X1 U348 ( .A(n754), .B(n755), .C(n756), .Y(n214) );
  INVX2 U349 ( .A(\CARRYB[11][9] ), .Y(n215) );
  INVX4 U350 ( .A(n215), .Y(n216) );
  AND2X1 U351 ( .A(n132), .B(n291), .Y(n952) );
  BUFX2 U352 ( .A(n578), .Y(n217) );
  BUFX2 U353 ( .A(n799), .Y(n218) );
  XNOR2X1 U354 ( .A(n220), .B(n444), .Y(\SUMB[10][5] ) );
  XOR2X1 U355 ( .A(\SUMB[11][4] ), .B(n222), .Y(n229) );
  XNOR2X1 U356 ( .A(n481), .B(n223), .Y(\SUMB[6][7] ) );
  INVX1 U357 ( .A(\SUMB[5][8] ), .Y(n223) );
  BUFX2 U358 ( .A(n800), .Y(n224) );
  XOR2X1 U359 ( .A(\CARRYB[9][6] ), .B(\ab[10][6] ), .Y(n228) );
  NAND2X1 U360 ( .A(\ab[14][2] ), .B(n389), .Y(n225) );
  INVX2 U361 ( .A(\SUMB[6][6] ), .Y(n308) );
  XNOR2X1 U362 ( .A(n226), .B(\SUMB[11][6] ), .Y(\SUMB[12][5] ) );
  XNOR2X1 U363 ( .A(\CARRYB[11][5] ), .B(\ab[12][5] ), .Y(n226) );
  XOR2X1 U364 ( .A(n227), .B(n89), .Y(\SUMB[15][1] ) );
  XOR2X1 U365 ( .A(\CARRYB[14][1] ), .B(\ab[15][1] ), .Y(n227) );
  XOR2X1 U366 ( .A(\SUMB[9][7] ), .B(n228), .Y(\SUMB[10][6] ) );
  XNOR2X1 U367 ( .A(n230), .B(\SUMB[13][6] ), .Y(\SUMB[14][5] ) );
  XNOR2X1 U368 ( .A(n97), .B(\ab[14][5] ), .Y(n230) );
  NAND3X1 U369 ( .A(n874), .B(n872), .C(n873), .Y(n231) );
  XOR2X1 U370 ( .A(n232), .B(n308), .Y(\SUMB[7][5] ) );
  XNOR2X1 U371 ( .A(\CARRYB[6][5] ), .B(\ab[7][5] ), .Y(n232) );
  XNOR2X1 U372 ( .A(n233), .B(\SUMB[9][11] ), .Y(\SUMB[10][10] ) );
  XNOR2X1 U373 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .Y(n233) );
  BUFX2 U374 ( .A(\SUMB[15][5] ), .Y(n234) );
  NAND3X1 U375 ( .A(n808), .B(n809), .C(n810), .Y(n235) );
  NAND3X1 U376 ( .A(n816), .B(n815), .C(n817), .Y(n236) );
  NAND3X1 U377 ( .A(n495), .B(n497), .C(n496), .Y(n237) );
  INVX2 U378 ( .A(\CARRYB[6][12] ), .Y(n238) );
  INVX4 U379 ( .A(n238), .Y(n239) );
  XOR2X1 U380 ( .A(n664), .B(n459), .Y(n240) );
  INVX2 U381 ( .A(\CARRYB[5][13] ), .Y(n241) );
  INVX4 U382 ( .A(n241), .Y(n242) );
  XOR2X1 U383 ( .A(n244), .B(n243), .Y(\SUMB[3][14] ) );
  XNOR2X1 U384 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .Y(n244) );
  NAND3X1 U385 ( .A(n472), .B(n471), .C(n473), .Y(n245) );
  AND2X2 U386 ( .A(n139), .B(\ab[0][14] ), .Y(n246) );
  XNOR2X1 U387 ( .A(n247), .B(n111), .Y(n852) );
  NAND3X1 U388 ( .A(n911), .B(n912), .C(n913), .Y(n249) );
  NAND2X1 U389 ( .A(\SUMB[4][6] ), .B(n56), .Y(n251) );
  NAND2X1 U390 ( .A(\SUMB[4][6] ), .B(\ab[5][5] ), .Y(n252) );
  NAND2X1 U391 ( .A(n56), .B(\ab[5][5] ), .Y(n253) );
  NAND3X1 U392 ( .A(n252), .B(n251), .C(n253), .Y(\CARRYB[5][5] ) );
  NAND2X1 U393 ( .A(n695), .B(n694), .Y(n254) );
  NAND3X1 U394 ( .A(n794), .B(n793), .C(n795), .Y(n255) );
  INVX1 U395 ( .A(n404), .Y(n256) );
  INVX2 U396 ( .A(\SUMB[2][12] ), .Y(n264) );
  XOR2X1 U397 ( .A(n51), .B(\ab[9][1] ), .Y(n257) );
  XOR2X1 U398 ( .A(n81), .B(n257), .Y(\SUMB[9][1] ) );
  NAND2X1 U399 ( .A(\SUMB[8][2] ), .B(\CARRYB[8][1] ), .Y(n258) );
  NAND2X1 U400 ( .A(\SUMB[8][2] ), .B(\ab[9][1] ), .Y(n259) );
  NAND2X1 U401 ( .A(\CARRYB[8][1] ), .B(\ab[9][1] ), .Y(n260) );
  NAND3X1 U402 ( .A(n259), .B(n258), .C(n260), .Y(\CARRYB[9][1] ) );
  NAND3X1 U403 ( .A(n724), .B(n722), .C(n723), .Y(n261) );
  XOR2X1 U404 ( .A(n53), .B(n262), .Y(\SUMB[7][1] ) );
  XOR2X1 U405 ( .A(\SUMB[6][2] ), .B(\ab[7][1] ), .Y(n262) );
  XNOR2X1 U406 ( .A(n975), .B(\ab[3][4] ), .Y(n624) );
  XOR2X1 U407 ( .A(n263), .B(n264), .Y(\SUMB[3][11] ) );
  XNOR2X1 U408 ( .A(\ab[3][11] ), .B(n165), .Y(n263) );
  AND2X1 U409 ( .A(n234), .B(\CARRYB[15][4] ), .Y(n956) );
  NAND2X1 U410 ( .A(\SUMB[10][6] ), .B(n255), .Y(n265) );
  NAND2X1 U411 ( .A(\SUMB[10][6] ), .B(\ab[11][5] ), .Y(n266) );
  NAND2X1 U412 ( .A(n255), .B(\ab[11][5] ), .Y(n267) );
  NAND3X1 U413 ( .A(n266), .B(n265), .C(n267), .Y(\CARRYB[11][5] ) );
  NAND3X1 U414 ( .A(n813), .B(n812), .C(n814), .Y(n268) );
  XNOR2X1 U415 ( .A(n269), .B(\SUMB[5][6] ), .Y(\SUMB[6][5] ) );
  XOR2X1 U416 ( .A(n662), .B(\ab[6][5] ), .Y(n269) );
  NAND3X1 U417 ( .A(n679), .B(n681), .C(n680), .Y(n270) );
  NAND3X1 U418 ( .A(n712), .B(n713), .C(n714), .Y(n271) );
  NAND3X1 U419 ( .A(n778), .B(n779), .C(n780), .Y(n272) );
  NAND3X1 U420 ( .A(n706), .B(n707), .C(n708), .Y(n273) );
  XNOR2X1 U421 ( .A(n274), .B(n6), .Y(\SUMB[9][7] ) );
  NAND2X1 U422 ( .A(\SUMB[11][4] ), .B(\CARRYB[11][3] ), .Y(n275) );
  NAND2X1 U423 ( .A(\CARRYB[11][3] ), .B(\ab[12][3] ), .Y(n276) );
  NAND2X1 U424 ( .A(\SUMB[11][4] ), .B(\ab[12][3] ), .Y(n277) );
  NAND3X1 U425 ( .A(n276), .B(n275), .C(n277), .Y(\CARRYB[12][3] ) );
  NAND3X1 U426 ( .A(n419), .B(n421), .C(n420), .Y(n278) );
  XOR2X1 U427 ( .A(\SUMB[4][11] ), .B(n279), .Y(n803) );
  XOR2X1 U428 ( .A(\CARRYB[7][8] ), .B(n280), .Y(n282) );
  XOR2X1 U429 ( .A(n281), .B(\SUMB[3][12] ), .Y(\SUMB[4][11] ) );
  XNOR2X1 U430 ( .A(n282), .B(n41), .Y(\SUMB[8][8] ) );
  XNOR2X1 U431 ( .A(n283), .B(\SUMB[4][9] ), .Y(\SUMB[5][8] ) );
  XOR2X1 U432 ( .A(\CARRYB[4][8] ), .B(n362), .Y(n283) );
  NAND3X1 U433 ( .A(n787), .B(n788), .C(n789), .Y(n284) );
  INVX2 U434 ( .A(\SUMB[9][6] ), .Y(n444) );
  INVX2 U435 ( .A(\CARRYB[5][12] ), .Y(n285) );
  INVX4 U436 ( .A(n285), .Y(n286) );
  XOR2X1 U437 ( .A(n287), .B(n106), .Y(\SUMB[4][8] ) );
  XOR2X1 U438 ( .A(\CARRYB[3][8] ), .B(\ab[4][8] ), .Y(n287) );
  XOR2X1 U439 ( .A(n288), .B(\SUMB[10][8] ), .Y(\SUMB[11][7] ) );
  XOR2X1 U440 ( .A(\CARRYB[10][7] ), .B(\ab[11][7] ), .Y(n288) );
  XNOR2X1 U441 ( .A(n290), .B(n289), .Y(\SUMB[8][9] ) );
  XOR2X1 U442 ( .A(\SUMB[7][10] ), .B(\ab[8][9] ), .Y(n290) );
  BUFX2 U443 ( .A(\SUMB[15][3] ), .Y(n291) );
  INVX1 U444 ( .A(\CARRYB[2][9] ), .Y(n875) );
  INVX1 U445 ( .A(n875), .Y(n876) );
  XNOR2X1 U446 ( .A(n292), .B(\SUMB[12][7] ), .Y(\SUMB[13][6] ) );
  XNOR2X1 U447 ( .A(\CARRYB[12][6] ), .B(\ab[13][6] ), .Y(n292) );
  XNOR2X1 U448 ( .A(\SUMB[15][5] ), .B(n293), .Y(\A1[18] ) );
  XNOR2X1 U449 ( .A(\ab[7][13] ), .B(n368), .Y(n629) );
  XNOR2X1 U450 ( .A(\SUMB[15][7] ), .B(n294), .Y(\A1[20] ) );
  XNOR2X1 U451 ( .A(\SUMB[3][13] ), .B(n295), .Y(\SUMB[4][12] ) );
  XNOR2X1 U452 ( .A(\CARRYB[3][12] ), .B(\ab[4][12] ), .Y(n295) );
  XNOR2X1 U453 ( .A(n629), .B(n296), .Y(\SUMB[7][13] ) );
  NAND2X1 U454 ( .A(\SUMB[4][7] ), .B(n284), .Y(n297) );
  NAND2X1 U455 ( .A(\SUMB[4][7] ), .B(\ab[5][6] ), .Y(n298) );
  NAND2X1 U456 ( .A(n284), .B(\ab[5][6] ), .Y(n299) );
  NAND3X1 U457 ( .A(n298), .B(n297), .C(n299), .Y(\CARRYB[5][6] ) );
  NAND3X1 U458 ( .A(n416), .B(n417), .C(n12), .Y(n300) );
  NAND3X1 U459 ( .A(n791), .B(n792), .C(n790), .Y(n301) );
  XOR2X1 U460 ( .A(n302), .B(\SUMB[14][1] ), .Y(\SUMB[15][0] ) );
  NAND2X1 U461 ( .A(n231), .B(\SUMB[14][1] ), .Y(n303) );
  NAND2X1 U462 ( .A(\SUMB[14][1] ), .B(\ab[15][0] ), .Y(n304) );
  NAND2X1 U463 ( .A(n231), .B(\ab[15][0] ), .Y(n305) );
  NAND3X1 U464 ( .A(n304), .B(n303), .C(n305), .Y(\CARRYB[15][0] ) );
  XNOR2X1 U465 ( .A(n306), .B(\SUMB[14][6] ), .Y(\SUMB[15][5] ) );
  XNOR2X1 U466 ( .A(\CARRYB[14][5] ), .B(\ab[15][5] ), .Y(n306) );
  XNOR2X1 U467 ( .A(n307), .B(\SUMB[5][9] ), .Y(\SUMB[6][8] ) );
  XNOR2X1 U468 ( .A(n372), .B(\SUMB[13][5] ), .Y(\SUMB[14][4] ) );
  XOR2X1 U469 ( .A(\CARRYB[9][3] ), .B(\ab[10][3] ), .Y(n314) );
  XOR2X1 U470 ( .A(\SUMB[3][3] ), .B(\ab[4][2] ), .Y(n309) );
  XOR2X1 U471 ( .A(n309), .B(n78), .Y(\SUMB[4][2] ) );
  NAND2X1 U472 ( .A(\CARRYB[3][2] ), .B(\SUMB[3][3] ), .Y(n310) );
  NAND2X1 U473 ( .A(\CARRYB[3][2] ), .B(\ab[4][2] ), .Y(n311) );
  NAND2X1 U474 ( .A(\SUMB[3][3] ), .B(\ab[4][2] ), .Y(n312) );
  NAND3X1 U475 ( .A(n311), .B(n310), .C(n312), .Y(\CARRYB[4][2] ) );
  BUFX2 U476 ( .A(\CARRYB[11][0] ), .Y(n313) );
  XNOR2X1 U477 ( .A(n314), .B(n425), .Y(\SUMB[10][3] ) );
  XOR2X1 U478 ( .A(n315), .B(n442), .Y(\SUMB[14][2] ) );
  XNOR2X1 U479 ( .A(n316), .B(n79), .Y(\SUMB[11][3] ) );
  XNOR2X1 U480 ( .A(\CARRYB[10][3] ), .B(\ab[11][3] ), .Y(n316) );
  NAND3X1 U481 ( .A(n583), .B(n584), .C(n585), .Y(n318) );
  XOR2X1 U482 ( .A(\CARRYB[2][6] ), .B(n319), .Y(n503) );
  NAND2X1 U483 ( .A(n1022), .B(n969), .Y(n319) );
  NAND2X1 U484 ( .A(\ab[12][1] ), .B(n982), .Y(n320) );
  BUFX2 U485 ( .A(\SUMB[4][3] ), .Y(n321) );
  BUFX2 U486 ( .A(\CARRYB[7][2] ), .Y(n322) );
  XOR2X1 U487 ( .A(n503), .B(n323), .Y(\SUMB[3][6] ) );
  INVX2 U488 ( .A(n1002), .Y(n905) );
  BUFX2 U489 ( .A(n688), .Y(n324) );
  NAND3X1 U490 ( .A(n599), .B(n598), .C(n597), .Y(n325) );
  XOR2X1 U491 ( .A(\CARRYB[14][6] ), .B(\ab[15][6] ), .Y(n326) );
  XOR2X1 U492 ( .A(\SUMB[14][7] ), .B(n326), .Y(\SUMB[15][6] ) );
  NAND2X1 U493 ( .A(\SUMB[14][7] ), .B(n11), .Y(n327) );
  NAND2X1 U494 ( .A(\SUMB[14][7] ), .B(\ab[15][6] ), .Y(n328) );
  NAND2X1 U495 ( .A(n11), .B(\ab[15][6] ), .Y(n329) );
  NAND3X1 U496 ( .A(n328), .B(n327), .C(n329), .Y(\CARRYB[15][6] ) );
  XOR2X1 U497 ( .A(\CARRYB[13][7] ), .B(\ab[14][7] ), .Y(n330) );
  XOR2X1 U498 ( .A(\SUMB[13][8] ), .B(n330), .Y(\SUMB[14][7] ) );
  NAND2X1 U499 ( .A(\SUMB[13][8] ), .B(\CARRYB[13][7] ), .Y(n331) );
  NAND2X1 U500 ( .A(\SUMB[13][8] ), .B(\ab[14][7] ), .Y(n332) );
  NAND2X1 U501 ( .A(\CARRYB[13][7] ), .B(\ab[14][7] ), .Y(n333) );
  NAND3X1 U502 ( .A(n332), .B(n331), .C(n333), .Y(\CARRYB[14][7] ) );
  INVX2 U503 ( .A(\CARRYB[6][7] ), .Y(n404) );
  NAND3X1 U504 ( .A(n925), .B(n926), .C(n927), .Y(n334) );
  NAND2X1 U505 ( .A(\ab[14][6] ), .B(n60), .Y(n335) );
  NAND2X1 U506 ( .A(\ab[14][6] ), .B(\SUMB[13][7] ), .Y(n336) );
  NAND2X1 U507 ( .A(n60), .B(\SUMB[13][7] ), .Y(n337) );
  NAND3X1 U508 ( .A(n335), .B(n336), .C(n337), .Y(\CARRYB[14][6] ) );
  NAND2X1 U509 ( .A(\ab[15][5] ), .B(n237), .Y(n338) );
  NAND2X1 U510 ( .A(\SUMB[14][6] ), .B(\ab[15][5] ), .Y(n339) );
  NAND2X1 U511 ( .A(n237), .B(n22), .Y(n340) );
  NAND3X1 U512 ( .A(n338), .B(n339), .C(n340), .Y(\CARRYB[15][5] ) );
  NAND2X1 U513 ( .A(n643), .B(n342), .Y(n343) );
  NAND2X1 U514 ( .A(n341), .B(\SUMB[12][8] ), .Y(n344) );
  NAND2X1 U515 ( .A(n343), .B(n344), .Y(\SUMB[13][7] ) );
  INVX1 U516 ( .A(n643), .Y(n341) );
  INVX1 U517 ( .A(\SUMB[12][8] ), .Y(n342) );
  NAND3X1 U518 ( .A(n853), .B(n854), .C(n855), .Y(n345) );
  NAND3X1 U519 ( .A(n908), .B(n909), .C(n910), .Y(n346) );
  INVX2 U520 ( .A(\SUMB[9][3] ), .Y(n347) );
  XOR2X1 U521 ( .A(\ab[2][2] ), .B(n960), .Y(n348) );
  XOR2X1 U522 ( .A(n348), .B(\SUMB[1][3] ), .Y(\SUMB[2][2] ) );
  XOR2X1 U523 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .Y(n349) );
  XOR2X1 U524 ( .A(n349), .B(n176), .Y(\SUMB[3][1] ) );
  NAND2X1 U525 ( .A(\ab[2][2] ), .B(n960), .Y(n350) );
  NAND2X1 U526 ( .A(\ab[2][2] ), .B(\SUMB[1][3] ), .Y(n351) );
  NAND2X1 U527 ( .A(n960), .B(\SUMB[1][3] ), .Y(n352) );
  NAND3X1 U528 ( .A(n350), .B(n351), .C(n352), .Y(\CARRYB[2][2] ) );
  NAND2X1 U529 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .Y(n353) );
  NAND2X1 U530 ( .A(\ab[3][1] ), .B(\SUMB[2][2] ), .Y(n354) );
  NAND2X1 U531 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n355) );
  NAND3X1 U532 ( .A(n353), .B(n354), .C(n355), .Y(\CARRYB[3][1] ) );
  XOR2X1 U533 ( .A(\SUMB[10][1] ), .B(\ab[11][0] ), .Y(n356) );
  XOR2X1 U534 ( .A(n967), .B(n356), .Y(\A1[9] ) );
  NAND2X1 U535 ( .A(n967), .B(\SUMB[10][1] ), .Y(n357) );
  NAND2X1 U536 ( .A(n967), .B(\ab[11][0] ), .Y(n358) );
  NAND2X1 U537 ( .A(\SUMB[10][1] ), .B(\ab[11][0] ), .Y(n359) );
  NAND3X1 U538 ( .A(n358), .B(n357), .C(n359), .Y(\CARRYB[11][0] ) );
  BUFX2 U539 ( .A(\SUMB[4][1] ), .Y(n360) );
  XNOR2X1 U540 ( .A(n361), .B(\SUMB[10][9] ), .Y(\SUMB[11][8] ) );
  XNOR2X1 U541 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .Y(n361) );
  XNOR2X1 U542 ( .A(n934), .B(n363), .Y(\SUMB[4][3] ) );
  INVX2 U543 ( .A(\SUMB[3][4] ), .Y(n363) );
  XOR2X1 U544 ( .A(n364), .B(n365), .Y(\SUMB[11][2] ) );
  XNOR2X1 U545 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .Y(n364) );
  INVX1 U546 ( .A(\SUMB[10][3] ), .Y(n365) );
  INVX2 U547 ( .A(\CARRYB[4][13] ), .Y(n366) );
  INVX4 U548 ( .A(n366), .Y(n367) );
  NAND3X1 U549 ( .A(n796), .B(n797), .C(n798), .Y(n369) );
  XOR2X1 U550 ( .A(n28), .B(n370), .Y(\SUMB[13][2] ) );
  XOR2X1 U551 ( .A(\CARRYB[12][2] ), .B(\ab[13][2] ), .Y(n370) );
  XOR2X1 U552 ( .A(n606), .B(n371), .Y(\SUMB[8][5] ) );
  INVX1 U553 ( .A(\SUMB[7][6] ), .Y(n371) );
  XNOR2X1 U554 ( .A(\CARRYB[13][4] ), .B(\ab[14][4] ), .Y(n372) );
  XOR2X1 U555 ( .A(n737), .B(n375), .Y(\SUMB[4][7] ) );
  INVX1 U556 ( .A(\SUMB[3][8] ), .Y(n375) );
  XNOR2X1 U557 ( .A(\ab[2][13] ), .B(n966), .Y(n914) );
  INVX2 U558 ( .A(n570), .Y(n571) );
  NAND3X1 U559 ( .A(n791), .B(n792), .C(n790), .Y(n376) );
  NAND3X1 U560 ( .A(n894), .B(n896), .C(n895), .Y(n377) );
  NAND2X1 U561 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(n378) );
  NAND2X1 U562 ( .A(\SUMB[7][4] ), .B(\ab[8][3] ), .Y(n379) );
  NAND2X1 U563 ( .A(\CARRYB[7][3] ), .B(\ab[8][3] ), .Y(n380) );
  NAND3X1 U564 ( .A(n379), .B(n378), .C(n380), .Y(\CARRYB[8][3] ) );
  XOR2X1 U565 ( .A(n906), .B(n381), .Y(n468) );
  NAND2X1 U566 ( .A(n59), .B(\SUMB[1][6] ), .Y(n382) );
  NAND2X1 U567 ( .A(n59), .B(\ab[2][5] ), .Y(n383) );
  NAND2X1 U568 ( .A(\SUMB[1][6] ), .B(\ab[2][5] ), .Y(n384) );
  NAND3X1 U569 ( .A(n383), .B(n382), .C(n384), .Y(\CARRYB[2][5] ) );
  AND2X2 U570 ( .A(B[7]), .B(A[2]), .Y(\ab[2][7] ) );
  NAND3X1 U571 ( .A(n889), .B(n890), .C(n888), .Y(n386) );
  NAND3X1 U572 ( .A(n945), .B(n946), .C(n947), .Y(n387) );
  NAND3X1 U573 ( .A(n553), .B(n551), .C(n552), .Y(n388) );
  NAND3X1 U574 ( .A(n920), .B(n921), .C(n919), .Y(n389) );
  NAND3X1 U575 ( .A(n893), .B(n892), .C(n891), .Y(n390) );
  NAND3X1 U576 ( .A(n801), .B(n218), .C(n224), .Y(n391) );
  NAND3X1 U577 ( .A(n687), .B(n324), .C(n689), .Y(n392) );
  NAND3X1 U578 ( .A(n862), .B(n91), .C(n863), .Y(n393) );
  NAND3X1 U579 ( .A(n901), .B(n902), .C(n161), .Y(n394) );
  NAND3X1 U580 ( .A(n842), .B(n843), .C(n844), .Y(n395) );
  NAND3X1 U581 ( .A(n556), .B(n554), .C(n555), .Y(n396) );
  NAND3X1 U582 ( .A(n922), .B(n923), .C(n924), .Y(n397) );
  NAND3X1 U583 ( .A(n768), .B(n769), .C(n770), .Y(n398) );
  BUFX2 U584 ( .A(n577), .Y(n399) );
  XNOR2X1 U585 ( .A(n705), .B(\ab[7][2] ), .Y(n449) );
  XNOR2X1 U586 ( .A(n837), .B(n400), .Y(\SUMB[13][1] ) );
  INVX2 U587 ( .A(n1016), .Y(n402) );
  INVX2 U588 ( .A(B[12]), .Y(n1010) );
  XOR2X1 U589 ( .A(n664), .B(n459), .Y(\SUMB[3][7] ) );
  NAND2X1 U590 ( .A(\ab[7][7] ), .B(n404), .Y(n405) );
  NAND2X1 U591 ( .A(n403), .B(n44), .Y(n406) );
  NAND2X1 U592 ( .A(n405), .B(n406), .Y(n897) );
  INVX1 U593 ( .A(\ab[7][7] ), .Y(n403) );
  NAND3X1 U594 ( .A(n587), .B(n588), .C(n589), .Y(n407) );
  XOR2X1 U595 ( .A(\SUMB[9][1] ), .B(\ab[10][0] ), .Y(n408) );
  XOR2X1 U596 ( .A(n52), .B(n408), .Y(\A1[8] ) );
  NAND2X1 U597 ( .A(\CARRYB[9][0] ), .B(\SUMB[9][1] ), .Y(n409) );
  NAND2X1 U598 ( .A(\CARRYB[9][0] ), .B(\ab[10][0] ), .Y(n410) );
  NAND2X1 U599 ( .A(\SUMB[9][1] ), .B(\ab[10][0] ), .Y(n411) );
  NAND3X1 U600 ( .A(n410), .B(n409), .C(n411), .Y(\CARRYB[10][0] ) );
  INVX1 U601 ( .A(\SUMB[7][2] ), .Y(n412) );
  INVX8 U602 ( .A(n1017), .Y(n1018) );
  XNOR2X1 U603 ( .A(n413), .B(\SUMB[2][4] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U604 ( .A(n983), .B(\ab[3][3] ), .Y(n413) );
  INVX2 U605 ( .A(n478), .Y(n414) );
  NOR2X1 U606 ( .A(n1017), .B(n1008), .Y(\ab[1][11] ) );
  XNOR2X1 U607 ( .A(n460), .B(n414), .Y(\SUMB[2][10] ) );
  AND2X2 U608 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(n415) );
  NAND2X1 U609 ( .A(\SUMB[5][7] ), .B(\ab[6][6] ), .Y(n416) );
  NAND2X1 U610 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .Y(n417) );
  NAND2X1 U611 ( .A(\SUMB[5][7] ), .B(\CARRYB[5][6] ), .Y(n418) );
  NAND3X1 U612 ( .A(n417), .B(n416), .C(n418), .Y(\CARRYB[6][6] ) );
  NAND2X1 U613 ( .A(\ab[7][5] ), .B(n334), .Y(n419) );
  NAND2X1 U614 ( .A(\SUMB[6][6] ), .B(\ab[7][5] ), .Y(n420) );
  NAND2X1 U615 ( .A(\SUMB[6][6] ), .B(n334), .Y(n421) );
  NAND3X1 U616 ( .A(n421), .B(n420), .C(n419), .Y(\CARRYB[7][5] ) );
  XNOR2X1 U617 ( .A(n422), .B(\SUMB[2][9] ), .Y(\SUMB[3][8] ) );
  XNOR2X1 U618 ( .A(n376), .B(n538), .Y(n422) );
  XOR2X1 U619 ( .A(n424), .B(\SUMB[6][5] ), .Y(\SUMB[7][4] ) );
  XOR2X1 U620 ( .A(\CARRYB[6][4] ), .B(\ab[7][4] ), .Y(n424) );
  INVX1 U621 ( .A(\SUMB[9][4] ), .Y(n425) );
  XOR2X1 U622 ( .A(\CARRYB[13][1] ), .B(\ab[14][1] ), .Y(n918) );
  XOR2X1 U623 ( .A(n48), .B(\ab[3][9] ), .Y(n596) );
  XOR2X1 U624 ( .A(\CARRYB[2][13] ), .B(\ab[3][13] ), .Y(n426) );
  XOR2X1 U625 ( .A(\SUMB[2][14] ), .B(n426), .Y(\SUMB[3][13] ) );
  NAND2X1 U626 ( .A(\SUMB[2][14] ), .B(n129), .Y(n427) );
  NAND2X1 U627 ( .A(\SUMB[2][14] ), .B(\ab[3][13] ), .Y(n428) );
  NAND2X1 U628 ( .A(n129), .B(\ab[3][13] ), .Y(n429) );
  NAND3X1 U629 ( .A(n428), .B(n427), .C(n429), .Y(\CARRYB[3][13] ) );
  XOR2X1 U630 ( .A(\ab[1][15] ), .B(\ab[2][14] ), .Y(n430) );
  XOR2X1 U631 ( .A(n430), .B(n30), .Y(\SUMB[2][14] ) );
  NAND2X1 U632 ( .A(n961), .B(\ab[1][15] ), .Y(n431) );
  NAND2X1 U633 ( .A(n961), .B(\ab[2][14] ), .Y(n432) );
  NAND2X1 U634 ( .A(\ab[1][15] ), .B(\ab[2][14] ), .Y(n433) );
  NAND3X1 U635 ( .A(n432), .B(n431), .C(n433), .Y(\CARRYB[2][14] ) );
  XOR2X1 U636 ( .A(\ab[2][11] ), .B(n506), .Y(n434) );
  XOR2X1 U637 ( .A(n434), .B(\SUMB[1][12] ), .Y(\SUMB[2][11] ) );
  XOR2X1 U638 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .Y(n435) );
  XOR2X1 U639 ( .A(n435), .B(\SUMB[2][11] ), .Y(\SUMB[3][10] ) );
  NAND2X1 U640 ( .A(\ab[2][11] ), .B(n506), .Y(n436) );
  NAND2X1 U641 ( .A(\ab[2][11] ), .B(\SUMB[1][12] ), .Y(n437) );
  NAND2X1 U642 ( .A(n506), .B(\SUMB[1][12] ), .Y(n438) );
  NAND3X1 U643 ( .A(n436), .B(n437), .C(n438), .Y(\CARRYB[2][11] ) );
  NAND2X1 U644 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .Y(n439) );
  NAND2X1 U645 ( .A(\ab[3][10] ), .B(\SUMB[2][11] ), .Y(n440) );
  NAND2X1 U646 ( .A(\CARRYB[2][10] ), .B(\SUMB[2][11] ), .Y(n441) );
  NAND3X1 U647 ( .A(n439), .B(n440), .C(n441), .Y(\CARRYB[3][10] ) );
  NAND3X1 U648 ( .A(n775), .B(n777), .C(n776), .Y(n443) );
  INVX2 U649 ( .A(\SUMB[7][7] ), .Y(n448) );
  BUFX2 U650 ( .A(\SUMB[1][5] ), .Y(n445) );
  BUFX2 U651 ( .A(\CARRYB[3][6] ), .Y(n446) );
  XOR2X1 U652 ( .A(n447), .B(n448), .Y(\SUMB[8][6] ) );
  XOR2X1 U653 ( .A(\SUMB[6][3] ), .B(n449), .Y(\SUMB[7][2] ) );
  NAND2X1 U654 ( .A(\SUMB[6][3] ), .B(\CARRYB[6][2] ), .Y(n450) );
  NAND2X1 U655 ( .A(\SUMB[6][3] ), .B(\ab[7][2] ), .Y(n451) );
  NAND2X1 U656 ( .A(\CARRYB[6][2] ), .B(\ab[7][2] ), .Y(n452) );
  NAND3X1 U657 ( .A(n451), .B(n450), .C(n452), .Y(\CARRYB[7][2] ) );
  XOR2X1 U658 ( .A(\CARRYB[8][2] ), .B(\ab[9][2] ), .Y(n453) );
  XOR2X1 U659 ( .A(n453), .B(n137), .Y(\SUMB[9][2] ) );
  NAND2X1 U660 ( .A(\SUMB[8][3] ), .B(n458), .Y(n454) );
  NAND2X1 U661 ( .A(\SUMB[8][3] ), .B(\ab[9][2] ), .Y(n455) );
  NAND2X1 U662 ( .A(n458), .B(\ab[9][2] ), .Y(n456) );
  NAND3X1 U663 ( .A(n455), .B(n454), .C(n456), .Y(\CARRYB[9][2] ) );
  NAND3X1 U664 ( .A(n532), .B(n533), .C(n534), .Y(n457) );
  NAND3X1 U665 ( .A(n565), .B(n564), .C(n566), .Y(n458) );
  INVX2 U666 ( .A(\SUMB[2][8] ), .Y(n459) );
  XOR2X1 U667 ( .A(\SUMB[1][11] ), .B(\ab[2][10] ), .Y(n460) );
  NAND2X1 U668 ( .A(\SUMB[1][11] ), .B(n478), .Y(n461) );
  NAND2X1 U669 ( .A(n478), .B(\ab[2][10] ), .Y(n462) );
  NAND2X1 U670 ( .A(\SUMB[1][11] ), .B(\ab[2][10] ), .Y(n463) );
  NAND3X1 U671 ( .A(n462), .B(n461), .C(n463), .Y(\CARRYB[2][10] ) );
  XNOR2X1 U672 ( .A(n395), .B(\ab[13][4] ), .Y(n464) );
  INVX1 U673 ( .A(\SUMB[1][10] ), .Y(n465) );
  NAND3X1 U674 ( .A(n898), .B(n899), .C(n900), .Y(n466) );
  NAND3X1 U675 ( .A(n579), .B(n581), .C(n580), .Y(n467) );
  XNOR2X1 U676 ( .A(n468), .B(\SUMB[1][8] ), .Y(\SUMB[2][7] ) );
  BUFX2 U677 ( .A(\SUMB[4][5] ), .Y(n469) );
  XOR2X1 U678 ( .A(\SUMB[1][7] ), .B(\ab[2][6] ), .Y(n470) );
  XOR2X1 U679 ( .A(n470), .B(n904), .Y(\SUMB[2][6] ) );
  NAND2X1 U680 ( .A(\SUMB[1][7] ), .B(n904), .Y(n471) );
  NAND2X1 U681 ( .A(n904), .B(\ab[2][6] ), .Y(n472) );
  NAND2X1 U682 ( .A(\SUMB[1][7] ), .B(\ab[2][6] ), .Y(n473) );
  NAND3X1 U683 ( .A(n472), .B(n471), .C(n473), .Y(\CARRYB[2][6] ) );
  NAND3X1 U684 ( .A(n225), .B(n486), .C(n487), .Y(n474) );
  NAND3X1 U685 ( .A(n784), .B(n785), .C(n786), .Y(n475) );
  XNOR2X1 U686 ( .A(\CARRYB[14][2] ), .B(n476), .Y(n686) );
  AND2X2 U687 ( .A(n181), .B(\ab[1][10] ), .Y(n478) );
  NAND3X1 U688 ( .A(n590), .B(n591), .C(n592), .Y(n479) );
  NAND3X1 U689 ( .A(n576), .B(n399), .C(n217), .Y(n480) );
  XOR2X1 U690 ( .A(n443), .B(\ab[6][7] ), .Y(n481) );
  NAND2X1 U691 ( .A(\SUMB[5][8] ), .B(\CARRYB[5][7] ), .Y(n482) );
  NAND2X1 U692 ( .A(\SUMB[5][8] ), .B(\ab[6][7] ), .Y(n483) );
  NAND2X1 U693 ( .A(\CARRYB[5][7] ), .B(\ab[6][7] ), .Y(n484) );
  NAND3X1 U694 ( .A(n483), .B(n482), .C(n484), .Y(\CARRYB[6][7] ) );
  NAND2X1 U695 ( .A(\ab[14][2] ), .B(n389), .Y(n485) );
  NAND2X1 U696 ( .A(\SUMB[13][3] ), .B(\ab[14][2] ), .Y(n486) );
  NAND2X1 U697 ( .A(\SUMB[13][3] ), .B(n389), .Y(n487) );
  NAND3X1 U698 ( .A(n485), .B(n486), .C(n487), .Y(\CARRYB[14][2] ) );
  NAND2X1 U699 ( .A(\ab[15][1] ), .B(n397), .Y(n488) );
  NAND2X1 U700 ( .A(\SUMB[14][2] ), .B(\ab[15][1] ), .Y(n489) );
  NAND2X1 U701 ( .A(\SUMB[14][2] ), .B(n397), .Y(n490) );
  NAND3X1 U702 ( .A(n488), .B(n490), .C(n489), .Y(\CARRYB[15][1] ) );
  INVX4 U703 ( .A(n997), .Y(n977) );
  INVX4 U704 ( .A(A[3]), .Y(n1021) );
  XNOR2X1 U705 ( .A(n491), .B(n75), .Y(\SUMB[5][3] ) );
  XNOR2X1 U706 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .Y(n491) );
  NAND2X1 U707 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .Y(n492) );
  NAND2X1 U708 ( .A(\SUMB[12][7] ), .B(\ab[13][6] ), .Y(n493) );
  NAND2X1 U709 ( .A(\CARRYB[12][6] ), .B(\SUMB[12][7] ), .Y(n494) );
  NAND3X1 U710 ( .A(n492), .B(n493), .C(n494), .Y(\CARRYB[13][6] ) );
  NAND2X1 U711 ( .A(\ab[14][5] ), .B(n97), .Y(n495) );
  NAND2X1 U712 ( .A(\SUMB[13][6] ), .B(\ab[14][5] ), .Y(n496) );
  NAND2X1 U713 ( .A(n97), .B(\SUMB[13][6] ), .Y(n497) );
  NAND3X1 U714 ( .A(n495), .B(n496), .C(n497), .Y(\CARRYB[14][5] ) );
  NAND2X1 U715 ( .A(\SUMB[10][8] ), .B(n235), .Y(n498) );
  NAND2X1 U716 ( .A(\SUMB[10][8] ), .B(\ab[11][7] ), .Y(n499) );
  NAND2X1 U717 ( .A(n235), .B(\ab[11][7] ), .Y(n500) );
  NAND3X1 U718 ( .A(n499), .B(n498), .C(n500), .Y(\CARRYB[11][7] ) );
  XNOR2X1 U719 ( .A(n387), .B(n501), .Y(n934) );
  NAND3X1 U720 ( .A(n859), .B(n860), .C(n861), .Y(n502) );
  XOR2X1 U721 ( .A(\CARRYB[12][4] ), .B(\ab[13][4] ), .Y(n811) );
  XNOR2X1 U722 ( .A(n504), .B(n254), .Y(\SUMB[14][3] ) );
  INVX1 U723 ( .A(n1051), .Y(n505) );
  INVX8 U724 ( .A(ZB), .Y(n1051) );
  AND2X2 U725 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(n506) );
  INVX1 U726 ( .A(n163), .Y(n1040) );
  BUFX4 U727 ( .A(B[9]), .Y(n507) );
  XOR2X1 U728 ( .A(n94), .B(\ab[6][4] ), .Y(n508) );
  NAND2X1 U729 ( .A(\SUMB[5][5] ), .B(\CARRYB[5][4] ), .Y(n509) );
  NAND2X1 U730 ( .A(\SUMB[5][5] ), .B(\ab[6][4] ), .Y(n510) );
  NAND2X1 U731 ( .A(\CARRYB[5][4] ), .B(\ab[6][4] ), .Y(n511) );
  NAND3X1 U732 ( .A(n511), .B(n510), .C(n509), .Y(\CARRYB[6][4] ) );
  XOR2X1 U733 ( .A(\CARRYB[9][9] ), .B(\ab[10][9] ), .Y(n512) );
  XOR2X1 U734 ( .A(\SUMB[9][10] ), .B(n512), .Y(\SUMB[10][9] ) );
  NAND2X1 U735 ( .A(\SUMB[9][10] ), .B(\CARRYB[9][9] ), .Y(n513) );
  NAND2X1 U736 ( .A(\SUMB[9][10] ), .B(\ab[10][9] ), .Y(n514) );
  NAND2X1 U737 ( .A(\CARRYB[9][9] ), .B(\ab[10][9] ), .Y(n515) );
  NAND3X1 U738 ( .A(n514), .B(n513), .C(n515), .Y(\CARRYB[10][9] ) );
  NAND2X1 U739 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .Y(n516) );
  NAND2X1 U740 ( .A(\ab[3][14] ), .B(\ab[2][15] ), .Y(n517) );
  NAND2X1 U741 ( .A(\CARRYB[2][14] ), .B(\ab[2][15] ), .Y(n518) );
  NAND3X1 U742 ( .A(n516), .B(n517), .C(n518), .Y(\CARRYB[3][14] ) );
  XOR2X1 U743 ( .A(\ab[4][14] ), .B(\ab[3][15] ), .Y(n519) );
  XOR2X1 U744 ( .A(n519), .B(\CARRYB[3][14] ), .Y(\SUMB[4][14] ) );
  NAND2X1 U745 ( .A(\ab[4][14] ), .B(\ab[3][15] ), .Y(n520) );
  NAND2X1 U746 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .Y(n521) );
  NAND2X1 U747 ( .A(\ab[3][15] ), .B(\CARRYB[3][14] ), .Y(n522) );
  NAND3X1 U748 ( .A(n520), .B(n521), .C(n522), .Y(\CARRYB[4][14] ) );
  NAND3X1 U749 ( .A(n749), .B(n750), .C(n751), .Y(n523) );
  NAND2X1 U750 ( .A(n527), .B(\CARRYB[3][1] ), .Y(n524) );
  NAND2X1 U751 ( .A(\ab[4][1] ), .B(n988), .Y(n525) );
  NAND2X1 U752 ( .A(n524), .B(n525), .Y(n616) );
  INVX1 U753 ( .A(\ab[4][1] ), .Y(n527) );
  INVX8 U754 ( .A(n1012), .Y(n1013) );
  INVX4 U755 ( .A(B[13]), .Y(n1012) );
  BUFX2 U756 ( .A(\SUMB[5][4] ), .Y(n526) );
  NAND3X1 U757 ( .A(n320), .B(n886), .C(n887), .Y(n528) );
  NAND3X1 U758 ( .A(n950), .B(n949), .C(n951), .Y(n529) );
  XNOR2X1 U759 ( .A(\ab[3][2] ), .B(n986), .Y(n730) );
  INVX2 U760 ( .A(n986), .Y(n987) );
  XNOR2X1 U761 ( .A(\CARRYB[4][9] ), .B(n530), .Y(n696) );
  BUFX2 U762 ( .A(A[0]), .Y(n531) );
  NAND2X1 U763 ( .A(\ab[5][3] ), .B(n180), .Y(n532) );
  NAND2X1 U764 ( .A(\ab[5][3] ), .B(\SUMB[4][4] ), .Y(n533) );
  NAND2X1 U765 ( .A(n180), .B(\SUMB[4][4] ), .Y(n534) );
  NAND3X1 U766 ( .A(n532), .B(n533), .C(n534), .Y(\CARRYB[5][3] ) );
  NAND2X1 U767 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .Y(n535) );
  NAND2X1 U768 ( .A(\ab[6][2] ), .B(\SUMB[5][3] ), .Y(n536) );
  NAND2X1 U769 ( .A(\CARRYB[5][2] ), .B(\SUMB[5][3] ), .Y(n537) );
  NAND3X1 U770 ( .A(n535), .B(n536), .C(n537), .Y(\CARRYB[6][2] ) );
  AND2X2 U771 ( .A(n1022), .B(n1005), .Y(n538) );
  INVX1 U772 ( .A(B[8]), .Y(n1004) );
  INVX4 U773 ( .A(n1004), .Y(n1005) );
  XOR2X1 U774 ( .A(\CARRYB[4][4] ), .B(\ab[5][4] ), .Y(n539) );
  XOR2X1 U775 ( .A(n469), .B(n539), .Y(\SUMB[5][4] ) );
  NAND2X1 U776 ( .A(\SUMB[4][5] ), .B(n479), .Y(n540) );
  NAND2X1 U777 ( .A(\SUMB[4][5] ), .B(\ab[5][4] ), .Y(n541) );
  NAND2X1 U778 ( .A(n479), .B(\ab[5][4] ), .Y(n542) );
  NAND3X1 U779 ( .A(n541), .B(n542), .C(n540), .Y(\CARRYB[5][4] ) );
  XNOR2X1 U780 ( .A(\ab[2][3] ), .B(n979), .Y(n729) );
  NAND3X1 U781 ( .A(n929), .B(n928), .C(n930), .Y(n543) );
  AND2X2 U782 ( .A(n984), .B(\ab[1][14] ), .Y(n961) );
  NAND3X1 U783 ( .A(n879), .B(n878), .C(n877), .Y(n544) );
  NAND2X1 U784 ( .A(\SUMB[7][2] ), .B(n261), .Y(n545) );
  NAND2X1 U785 ( .A(\SUMB[7][2] ), .B(\ab[8][1] ), .Y(n546) );
  NAND2X1 U786 ( .A(n261), .B(\ab[8][1] ), .Y(n547) );
  NAND3X1 U787 ( .A(n546), .B(n545), .C(n547), .Y(\CARRYB[8][1] ) );
  BUFX2 U788 ( .A(\SUMB[12][1] ), .Y(n548) );
  NAND3X1 U789 ( .A(n626), .B(n625), .C(n627), .Y(n549) );
  XOR2X1 U790 ( .A(\SUMB[11][1] ), .B(\ab[12][0] ), .Y(n550) );
  XOR2X1 U791 ( .A(n313), .B(n550), .Y(\A1[10] ) );
  NAND2X1 U792 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Y(n551) );
  NAND2X1 U793 ( .A(\CARRYB[11][0] ), .B(\ab[12][0] ), .Y(n552) );
  NAND2X1 U794 ( .A(\SUMB[11][1] ), .B(\ab[12][0] ), .Y(n553) );
  NAND3X1 U795 ( .A(n553), .B(n552), .C(n551), .Y(\CARRYB[12][0] ) );
  NAND2X1 U796 ( .A(\ab[2][7] ), .B(n73), .Y(n554) );
  NAND2X1 U797 ( .A(\SUMB[1][8] ), .B(n73), .Y(n555) );
  NAND2X1 U798 ( .A(\SUMB[1][8] ), .B(\ab[2][7] ), .Y(n556) );
  NAND3X1 U799 ( .A(n556), .B(n555), .C(n554), .Y(\CARRYB[2][7] ) );
  NAND2X1 U800 ( .A(\ab[3][6] ), .B(n245), .Y(n557) );
  NAND2X1 U801 ( .A(\SUMB[2][7] ), .B(\ab[3][6] ), .Y(n558) );
  NAND2X1 U802 ( .A(\SUMB[2][7] ), .B(n245), .Y(n559) );
  NAND3X1 U803 ( .A(n557), .B(n558), .C(n559), .Y(\CARRYB[3][6] ) );
  NAND2X1 U804 ( .A(\SUMB[1][10] ), .B(\ab[2][9] ), .Y(n560) );
  NAND2X1 U805 ( .A(\SUMB[1][10] ), .B(n760), .Y(n561) );
  NAND2X1 U806 ( .A(n760), .B(\ab[2][9] ), .Y(n562) );
  NAND3X1 U807 ( .A(n561), .B(n560), .C(n562), .Y(\CARRYB[2][9] ) );
  XNOR2X1 U808 ( .A(n569), .B(\SUMB[9][9] ), .Y(\SUMB[10][8] ) );
  XOR2X1 U809 ( .A(\SUMB[7][3] ), .B(\ab[8][2] ), .Y(n563) );
  XOR2X1 U810 ( .A(n322), .B(n563), .Y(\SUMB[8][2] ) );
  NAND2X1 U811 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(n564) );
  NAND2X1 U812 ( .A(\CARRYB[7][2] ), .B(\ab[8][2] ), .Y(n565) );
  NAND2X1 U813 ( .A(\SUMB[7][3] ), .B(\ab[8][2] ), .Y(n566) );
  NAND3X1 U814 ( .A(n565), .B(n564), .C(n566), .Y(\CARRYB[8][2] ) );
  XNOR2X1 U815 ( .A(n567), .B(n445), .Y(\SUMB[2][4] ) );
  XNOR2X1 U816 ( .A(n654), .B(\ab[2][4] ), .Y(n567) );
  AND2X2 U817 ( .A(n4), .B(n1015), .Y(\ab[2][14] ) );
  XOR2X1 U818 ( .A(n568), .B(n570), .Y(n745) );
  XNOR2X1 U819 ( .A(\CARRYB[9][8] ), .B(\ab[10][8] ), .Y(n569) );
  INVX2 U820 ( .A(\CARRYB[11][7] ), .Y(n570) );
  NAND2X1 U821 ( .A(\SUMB[3][6] ), .B(\CARRYB[3][5] ), .Y(n572) );
  NAND2X1 U822 ( .A(\SUMB[3][6] ), .B(\ab[4][5] ), .Y(n573) );
  NAND2X1 U823 ( .A(\CARRYB[3][5] ), .B(\ab[4][5] ), .Y(n574) );
  NAND3X1 U824 ( .A(n574), .B(n572), .C(n573), .Y(\CARRYB[4][5] ) );
  XOR2X1 U825 ( .A(n575), .B(\SUMB[7][8] ), .Y(\SUMB[8][7] ) );
  NAND2X1 U826 ( .A(\ab[7][8] ), .B(n466), .Y(n576) );
  NAND2X1 U827 ( .A(\SUMB[6][9] ), .B(\ab[7][8] ), .Y(n577) );
  NAND2X1 U828 ( .A(n466), .B(\SUMB[6][9] ), .Y(n578) );
  NAND3X1 U829 ( .A(n576), .B(n577), .C(n578), .Y(\CARRYB[7][8] ) );
  NAND2X1 U830 ( .A(\ab[8][7] ), .B(n394), .Y(n579) );
  NAND2X1 U831 ( .A(\SUMB[7][8] ), .B(\ab[8][7] ), .Y(n580) );
  NAND2X1 U832 ( .A(\SUMB[7][8] ), .B(n394), .Y(n581) );
  NAND3X1 U833 ( .A(n579), .B(n580), .C(n581), .Y(\CARRYB[8][7] ) );
  NAND3X1 U834 ( .A(n715), .B(n717), .C(n716), .Y(n582) );
  NAND2X1 U835 ( .A(\SUMB[6][7] ), .B(n300), .Y(n583) );
  NAND2X1 U836 ( .A(\SUMB[6][7] ), .B(\ab[7][6] ), .Y(n584) );
  NAND2X1 U837 ( .A(n300), .B(\ab[7][6] ), .Y(n585) );
  NAND3X1 U838 ( .A(n585), .B(n583), .C(n584), .Y(\CARRYB[7][6] ) );
  INVX1 U839 ( .A(n1013), .Y(n1038) );
  INVX2 U840 ( .A(n981), .Y(n982) );
  NOR2X1 U841 ( .A(n1012), .B(n655), .Y(\ab[0][13] ) );
  XOR2X1 U842 ( .A(\CARRYB[3][4] ), .B(\ab[4][4] ), .Y(n586) );
  XOR2X1 U843 ( .A(\SUMB[3][5] ), .B(n586), .Y(\SUMB[4][4] ) );
  NAND2X1 U844 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .Y(n587) );
  NAND2X1 U845 ( .A(\SUMB[2][6] ), .B(\ab[3][5] ), .Y(n588) );
  NAND2X1 U846 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n589) );
  NAND3X1 U847 ( .A(n587), .B(n588), .C(n589), .Y(\CARRYB[3][5] ) );
  NAND2X1 U848 ( .A(\ab[4][4] ), .B(n549), .Y(n590) );
  NAND2X1 U849 ( .A(\SUMB[3][5] ), .B(\ab[4][4] ), .Y(n591) );
  NAND2X1 U850 ( .A(\SUMB[3][5] ), .B(n549), .Y(n592) );
  NAND3X1 U851 ( .A(n590), .B(n591), .C(n592), .Y(\CARRYB[4][4] ) );
  INVX1 U852 ( .A(n662), .Y(n663) );
  XNOR2X1 U853 ( .A(n803), .B(n112), .Y(\SUMB[5][10] ) );
  XNOR2X1 U854 ( .A(n594), .B(\SUMB[1][13] ), .Y(\SUMB[2][12] ) );
  XNOR2X1 U855 ( .A(n802), .B(\ab[2][12] ), .Y(n594) );
  XNOR2X1 U856 ( .A(n595), .B(\SUMB[14][4] ), .Y(\SUMB[15][3] ) );
  XOR2X1 U857 ( .A(n219), .B(n596), .Y(\SUMB[3][9] ) );
  NAND2X1 U858 ( .A(\SUMB[2][10] ), .B(n876), .Y(n597) );
  NAND2X1 U859 ( .A(\SUMB[2][10] ), .B(\ab[3][9] ), .Y(n598) );
  NAND2X1 U860 ( .A(n876), .B(\ab[3][9] ), .Y(n599) );
  NAND3X1 U861 ( .A(n598), .B(n597), .C(n599), .Y(\CARRYB[3][9] ) );
  NAND3X1 U862 ( .A(n882), .B(n881), .C(n880), .Y(n600) );
  NAND3X1 U863 ( .A(n772), .B(n773), .C(n774), .Y(n601) );
  XOR2X1 U864 ( .A(\CARRYB[8][4] ), .B(\ab[9][4] ), .Y(n602) );
  XOR2X1 U865 ( .A(\SUMB[8][5] ), .B(n602), .Y(\SUMB[9][4] ) );
  NAND2X1 U866 ( .A(\SUMB[8][5] ), .B(n544), .Y(n603) );
  NAND2X1 U867 ( .A(\SUMB[8][5] ), .B(\ab[9][4] ), .Y(n604) );
  NAND2X1 U868 ( .A(n544), .B(\ab[9][4] ), .Y(n605) );
  NAND3X1 U869 ( .A(n605), .B(n604), .C(n603), .Y(\CARRYB[9][4] ) );
  XNOR2X1 U870 ( .A(\CARRYB[7][5] ), .B(\ab[8][5] ), .Y(n606) );
  BUFX2 U871 ( .A(\SUMB[15][0] ), .Y(n607) );
  XOR2X1 U872 ( .A(n86), .B(\ab[8][0] ), .Y(n608) );
  XOR2X1 U873 ( .A(n608), .B(n85), .Y(\A1[6] ) );
  NAND2X1 U874 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(n609) );
  NAND2X1 U875 ( .A(\CARRYB[7][0] ), .B(\ab[8][0] ), .Y(n610) );
  NAND2X1 U876 ( .A(\SUMB[7][1] ), .B(\ab[8][0] ), .Y(n611) );
  NAND3X1 U877 ( .A(n611), .B(n609), .C(n610), .Y(\CARRYB[8][0] ) );
  XOR2X1 U878 ( .A(\SUMB[6][1] ), .B(\ab[7][0] ), .Y(n612) );
  XOR2X1 U879 ( .A(\CARRYB[6][0] ), .B(n612), .Y(\A1[5] ) );
  NAND2X1 U880 ( .A(\CARRYB[6][0] ), .B(\SUMB[6][1] ), .Y(n613) );
  NAND2X1 U881 ( .A(\CARRYB[6][0] ), .B(\ab[7][0] ), .Y(n614) );
  NAND2X1 U882 ( .A(\SUMB[6][1] ), .B(\ab[7][0] ), .Y(n615) );
  NAND3X1 U883 ( .A(n615), .B(n613), .C(n614), .Y(\CARRYB[7][0] ) );
  XOR2X1 U884 ( .A(n616), .B(\SUMB[3][2] ), .Y(\SUMB[4][1] ) );
  XOR2X1 U885 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .Y(n617) );
  XOR2X1 U886 ( .A(n617), .B(n360), .Y(\A1[3] ) );
  NAND2X1 U887 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .Y(n618) );
  NAND2X1 U888 ( .A(\ab[4][1] ), .B(\SUMB[3][2] ), .Y(n619) );
  NAND2X1 U889 ( .A(\CARRYB[3][1] ), .B(\SUMB[3][2] ), .Y(n620) );
  NAND3X1 U890 ( .A(n618), .B(n619), .C(n620), .Y(\CARRYB[4][1] ) );
  NAND2X1 U891 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .Y(n621) );
  NAND2X1 U892 ( .A(\ab[5][0] ), .B(\SUMB[4][1] ), .Y(n622) );
  NAND2X1 U893 ( .A(\CARRYB[4][0] ), .B(\SUMB[4][1] ), .Y(n623) );
  NAND3X1 U894 ( .A(n621), .B(n622), .C(n623), .Y(\CARRYB[5][0] ) );
  XOR2X1 U895 ( .A(n98), .B(n624), .Y(\SUMB[3][4] ) );
  NAND2X1 U896 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n625) );
  NAND2X1 U897 ( .A(\SUMB[2][5] ), .B(\ab[3][4] ), .Y(n626) );
  NAND2X1 U898 ( .A(\CARRYB[2][4] ), .B(\ab[3][4] ), .Y(n627) );
  NAND3X1 U899 ( .A(n626), .B(n625), .C(n627), .Y(\CARRYB[3][4] ) );
  XOR2X1 U900 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .Y(n628) );
  XOR2X1 U901 ( .A(n628), .B(\ab[5][15] ), .Y(\SUMB[6][14] ) );
  NAND2X1 U902 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .Y(n630) );
  NAND2X1 U903 ( .A(\ab[6][14] ), .B(\ab[5][15] ), .Y(n631) );
  NAND2X1 U904 ( .A(\CARRYB[5][14] ), .B(\ab[5][15] ), .Y(n632) );
  NAND3X1 U905 ( .A(n630), .B(n631), .C(n632), .Y(\CARRYB[6][14] ) );
  NAND2X1 U906 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .Y(n633) );
  NAND2X1 U907 ( .A(\ab[7][13] ), .B(\SUMB[6][14] ), .Y(n634) );
  NAND2X1 U908 ( .A(\CARRYB[6][13] ), .B(\SUMB[6][14] ), .Y(n635) );
  NAND3X1 U909 ( .A(n633), .B(n634), .C(n635), .Y(\CARRYB[7][13] ) );
  NAND2X1 U910 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .Y(n636) );
  NAND2X1 U911 ( .A(\SUMB[8][12] ), .B(\ab[9][11] ), .Y(n637) );
  NAND2X1 U912 ( .A(\CARRYB[8][11] ), .B(\SUMB[8][12] ), .Y(n638) );
  NAND3X1 U913 ( .A(n636), .B(n637), .C(n638), .Y(\CARRYB[9][11] ) );
  NAND2X1 U914 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .Y(n639) );
  NAND2X1 U915 ( .A(\SUMB[9][11] ), .B(\ab[10][10] ), .Y(n640) );
  NAND2X1 U916 ( .A(\CARRYB[9][10] ), .B(\SUMB[9][11] ), .Y(n641) );
  NAND3X1 U917 ( .A(n639), .B(n640), .C(n641), .Y(\CARRYB[10][10] ) );
  XOR2X1 U918 ( .A(n642), .B(\SUMB[11][9] ), .Y(\SUMB[12][8] ) );
  XOR2X1 U919 ( .A(\CARRYB[12][7] ), .B(\ab[13][7] ), .Y(n643) );
  NAND2X1 U920 ( .A(\ab[12][8] ), .B(n20), .Y(n644) );
  NAND2X1 U921 ( .A(\ab[12][8] ), .B(\SUMB[11][9] ), .Y(n645) );
  NAND2X1 U922 ( .A(n20), .B(\SUMB[11][9] ), .Y(n646) );
  NAND3X1 U923 ( .A(n644), .B(n645), .C(n646), .Y(\CARRYB[12][8] ) );
  NAND2X1 U924 ( .A(\ab[13][7] ), .B(n523), .Y(n647) );
  NAND2X1 U925 ( .A(\ab[13][7] ), .B(\SUMB[12][8] ), .Y(n648) );
  NAND2X1 U926 ( .A(n523), .B(\SUMB[12][8] ), .Y(n649) );
  NAND3X1 U927 ( .A(n647), .B(n648), .C(n649), .Y(\CARRYB[13][7] ) );
  XOR2X1 U928 ( .A(\CARRYB[7][12] ), .B(\ab[8][12] ), .Y(n650) );
  XOR2X1 U929 ( .A(\SUMB[7][13] ), .B(n650), .Y(\SUMB[8][12] ) );
  NAND2X1 U930 ( .A(\SUMB[7][13] ), .B(n214), .Y(n651) );
  NAND2X1 U931 ( .A(\SUMB[7][13] ), .B(\ab[8][12] ), .Y(n652) );
  NAND2X1 U932 ( .A(n214), .B(\ab[8][12] ), .Y(n653) );
  NAND3X1 U933 ( .A(n652), .B(n651), .C(n653), .Y(\CARRYB[8][12] ) );
  AND2X2 U934 ( .A(n962), .B(\ab[1][4] ), .Y(n654) );
  INVX2 U935 ( .A(n907), .Y(n984) );
  NAND2X1 U936 ( .A(n49), .B(\ab[10][3] ), .Y(n656) );
  NAND2X1 U937 ( .A(\SUMB[9][4] ), .B(n49), .Y(n657) );
  NAND2X1 U938 ( .A(\ab[10][3] ), .B(\SUMB[9][4] ), .Y(n658) );
  NAND3X1 U939 ( .A(n656), .B(n657), .C(n658), .Y(\CARRYB[10][3] ) );
  NAND2X1 U940 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .Y(n659) );
  NAND2X1 U941 ( .A(\ab[11][2] ), .B(\SUMB[10][3] ), .Y(n660) );
  NAND2X1 U942 ( .A(\SUMB[10][3] ), .B(\CARRYB[10][2] ), .Y(n661) );
  NAND3X1 U943 ( .A(n659), .B(n660), .C(n661), .Y(\CARRYB[11][2] ) );
  INVX2 U944 ( .A(\CARRYB[5][5] ), .Y(n662) );
  XNOR2X1 U945 ( .A(\CARRYB[2][7] ), .B(\ab[3][7] ), .Y(n664) );
  XOR2X1 U946 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .Y(n665) );
  XOR2X1 U947 ( .A(n665), .B(\SUMB[7][11] ), .Y(\SUMB[8][10] ) );
  NAND2X1 U948 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .Y(n666) );
  NAND2X1 U949 ( .A(\ab[7][11] ), .B(\SUMB[6][12] ), .Y(n667) );
  NAND2X1 U950 ( .A(\CARRYB[6][11] ), .B(\SUMB[6][12] ), .Y(n668) );
  NAND3X1 U951 ( .A(n666), .B(n667), .C(n668), .Y(\CARRYB[7][11] ) );
  NAND2X1 U952 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .Y(n669) );
  NAND2X1 U953 ( .A(\ab[8][10] ), .B(\SUMB[7][11] ), .Y(n670) );
  NAND2X1 U954 ( .A(\CARRYB[7][10] ), .B(\SUMB[7][11] ), .Y(n671) );
  NAND3X1 U955 ( .A(n669), .B(n670), .C(n671), .Y(\CARRYB[8][10] ) );
  XOR2X1 U956 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .Y(n672) );
  XOR2X1 U957 ( .A(n672), .B(\SUMB[8][10] ), .Y(\SUMB[9][9] ) );
  NAND2X1 U958 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .Y(n673) );
  NAND2X1 U959 ( .A(\ab[9][9] ), .B(\SUMB[8][10] ), .Y(n674) );
  NAND2X1 U960 ( .A(\CARRYB[8][9] ), .B(\SUMB[8][10] ), .Y(n675) );
  NAND3X1 U961 ( .A(n673), .B(n674), .C(n675), .Y(\CARRYB[9][9] ) );
  NAND2X1 U962 ( .A(\ab[10][8] ), .B(n55), .Y(n676) );
  NAND2X1 U963 ( .A(\ab[10][8] ), .B(\SUMB[9][9] ), .Y(n677) );
  NAND2X1 U964 ( .A(n55), .B(\SUMB[9][9] ), .Y(n678) );
  NAND3X1 U965 ( .A(n676), .B(n677), .C(n678), .Y(\CARRYB[10][8] ) );
  NAND2X1 U966 ( .A(\ab[14][4] ), .B(n268), .Y(n679) );
  NAND2X1 U967 ( .A(\SUMB[13][5] ), .B(\ab[14][4] ), .Y(n680) );
  NAND2X1 U968 ( .A(\SUMB[13][5] ), .B(n268), .Y(n681) );
  NAND3X1 U969 ( .A(n679), .B(n680), .C(n681), .Y(\CARRYB[14][4] ) );
  NAND2X1 U970 ( .A(\ab[15][3] ), .B(n392), .Y(n682) );
  NAND2X1 U971 ( .A(\SUMB[14][4] ), .B(\ab[15][3] ), .Y(n683) );
  NAND2X1 U972 ( .A(\SUMB[14][4] ), .B(n392), .Y(n684) );
  NAND3X1 U973 ( .A(n682), .B(n683), .C(n684), .Y(\CARRYB[15][3] ) );
  XNOR2X1 U974 ( .A(n685), .B(\SUMB[11][7] ), .Y(\SUMB[12][6] ) );
  XNOR2X1 U975 ( .A(\CARRYB[11][6] ), .B(\ab[12][6] ), .Y(n685) );
  XOR2X1 U976 ( .A(n686), .B(n133), .Y(\SUMB[15][2] ) );
  NAND2X1 U977 ( .A(\ab[14][3] ), .B(n134), .Y(n687) );
  NAND2X1 U978 ( .A(\ab[14][3] ), .B(\SUMB[13][4] ), .Y(n688) );
  NAND2X1 U979 ( .A(n134), .B(\SUMB[13][4] ), .Y(n689) );
  NAND3X1 U980 ( .A(n687), .B(n688), .C(n689), .Y(\CARRYB[14][3] ) );
  NAND2X1 U981 ( .A(\ab[15][2] ), .B(n474), .Y(n690) );
  NAND2X1 U982 ( .A(\ab[15][2] ), .B(\SUMB[14][3] ), .Y(n691) );
  NAND2X1 U983 ( .A(n474), .B(\SUMB[14][3] ), .Y(n692) );
  NAND3X1 U984 ( .A(n690), .B(n692), .C(n691), .Y(\CARRYB[15][2] ) );
  NAND2X1 U985 ( .A(\SUMB[12][5] ), .B(n464), .Y(n694) );
  NAND2X1 U986 ( .A(n693), .B(n811), .Y(n695) );
  NAND2X1 U987 ( .A(n695), .B(n694), .Y(\SUMB[13][4] ) );
  INVX1 U988 ( .A(\SUMB[12][5] ), .Y(n693) );
  XOR2X1 U989 ( .A(n696), .B(\SUMB[4][10] ), .Y(\SUMB[5][9] ) );
  NAND2X1 U990 ( .A(\ab[5][9] ), .B(n502), .Y(n697) );
  NAND2X1 U991 ( .A(\ab[5][9] ), .B(\SUMB[4][10] ), .Y(n698) );
  NAND2X1 U992 ( .A(\SUMB[4][10] ), .B(n502), .Y(n699) );
  NAND3X1 U993 ( .A(n697), .B(n698), .C(n699), .Y(\CARRYB[5][9] ) );
  NAND2X1 U994 ( .A(\SUMB[5][10] ), .B(\ab[6][9] ), .Y(n700) );
  NAND2X1 U995 ( .A(\CARRYB[5][9] ), .B(\ab[6][9] ), .Y(n701) );
  NAND2X1 U996 ( .A(\SUMB[5][10] ), .B(\CARRYB[5][9] ), .Y(n702) );
  NAND3X1 U997 ( .A(n700), .B(n701), .C(n702), .Y(\CARRYB[6][9] ) );
  NAND3X1 U998 ( .A(n842), .B(n843), .C(n844), .Y(n703) );
  BUFX2 U999 ( .A(\SUMB[13][1] ), .Y(n704) );
  AND2X2 U1000 ( .A(\SUMB[15][1] ), .B(\CARRYB[15][0] ), .Y(n955) );
  INVX2 U1001 ( .A(\CARRYB[6][2] ), .Y(n705) );
  NAND2X1 U1002 ( .A(\ab[11][6] ), .B(n88), .Y(n706) );
  NAND2X1 U1003 ( .A(\SUMB[10][7] ), .B(\ab[11][6] ), .Y(n707) );
  NAND2X1 U1004 ( .A(\SUMB[10][7] ), .B(n88), .Y(n708) );
  NAND3X1 U1005 ( .A(n706), .B(n707), .C(n708), .Y(\CARRYB[11][6] ) );
  NAND2X1 U1006 ( .A(\ab[12][5] ), .B(n154), .Y(n709) );
  NAND2X1 U1007 ( .A(\SUMB[11][6] ), .B(\ab[12][5] ), .Y(n710) );
  NAND2X1 U1008 ( .A(n154), .B(\SUMB[11][6] ), .Y(n711) );
  NAND3X1 U1009 ( .A(n709), .B(n710), .C(n711), .Y(\CARRYB[12][5] ) );
  NAND2X1 U1010 ( .A(n160), .B(n183), .Y(n712) );
  NAND2X1 U1011 ( .A(\SUMB[1][13] ), .B(n183), .Y(n713) );
  NAND2X1 U1012 ( .A(\SUMB[1][13] ), .B(n160), .Y(n714) );
  NAND3X1 U1013 ( .A(n712), .B(n713), .C(n714), .Y(\CARRYB[2][12] ) );
  NAND2X1 U1014 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .Y(n715) );
  NAND2X1 U1015 ( .A(\SUMB[2][12] ), .B(\ab[3][11] ), .Y(n716) );
  NAND2X1 U1016 ( .A(\SUMB[2][12] ), .B(\CARRYB[2][11] ), .Y(n717) );
  NAND3X1 U1017 ( .A(n715), .B(n716), .C(n717), .Y(\CARRYB[3][11] ) );
  XNOR2X1 U1018 ( .A(n718), .B(\SUMB[9][8] ), .Y(\SUMB[10][7] ) );
  XNOR2X1 U1019 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .Y(n718) );
  NAND2X1 U1020 ( .A(n7), .B(\SUMB[9][2] ), .Y(n719) );
  NAND2X1 U1021 ( .A(\CARRYB[9][1] ), .B(\ab[10][1] ), .Y(n720) );
  NAND2X1 U1022 ( .A(\SUMB[9][2] ), .B(\ab[10][1] ), .Y(n721) );
  NAND3X1 U1023 ( .A(n720), .B(n721), .C(n719), .Y(\CARRYB[10][1] ) );
  NAND2X1 U1024 ( .A(\SUMB[6][2] ), .B(\CARRYB[6][1] ), .Y(n722) );
  NAND2X1 U1025 ( .A(\CARRYB[6][1] ), .B(\ab[7][1] ), .Y(n723) );
  NAND2X1 U1026 ( .A(\SUMB[6][2] ), .B(\ab[7][1] ), .Y(n724) );
  NAND3X1 U1027 ( .A(n724), .B(n722), .C(n723), .Y(\CARRYB[7][1] ) );
  XOR2X1 U1028 ( .A(\CARRYB[4][1] ), .B(\ab[5][1] ), .Y(n725) );
  XOR2X1 U1029 ( .A(\SUMB[4][2] ), .B(n725), .Y(\SUMB[5][1] ) );
  NAND2X1 U1030 ( .A(\SUMB[4][2] ), .B(\CARRYB[4][1] ), .Y(n726) );
  NAND2X1 U1031 ( .A(\SUMB[4][2] ), .B(\ab[5][1] ), .Y(n727) );
  NAND2X1 U1032 ( .A(\CARRYB[4][1] ), .B(\ab[5][1] ), .Y(n728) );
  NAND3X1 U1033 ( .A(n727), .B(n728), .C(n726), .Y(\CARRYB[5][1] ) );
  XOR2X1 U1034 ( .A(n729), .B(\SUMB[1][4] ), .Y(\SUMB[2][3] ) );
  XOR2X1 U1035 ( .A(n730), .B(\SUMB[2][3] ), .Y(\SUMB[3][2] ) );
  NAND2X1 U1036 ( .A(\ab[2][3] ), .B(n959), .Y(n731) );
  NAND2X1 U1037 ( .A(\ab[2][3] ), .B(\SUMB[1][4] ), .Y(n732) );
  NAND2X1 U1038 ( .A(n959), .B(\SUMB[1][4] ), .Y(n733) );
  NAND3X1 U1039 ( .A(n731), .B(n732), .C(n733), .Y(\CARRYB[2][3] ) );
  NAND2X1 U1040 ( .A(\ab[3][2] ), .B(n987), .Y(n734) );
  NAND2X1 U1041 ( .A(\ab[3][2] ), .B(\SUMB[2][3] ), .Y(n735) );
  NAND2X1 U1042 ( .A(n987), .B(\SUMB[2][3] ), .Y(n736) );
  NAND3X1 U1043 ( .A(n734), .B(n735), .C(n736), .Y(\CARRYB[3][2] ) );
  XNOR2X1 U1044 ( .A(\CARRYB[3][7] ), .B(\ab[4][7] ), .Y(n737) );
  NAND2X1 U1045 ( .A(\SUMB[6][4] ), .B(n529), .Y(n738) );
  NAND2X1 U1046 ( .A(\SUMB[6][4] ), .B(\ab[7][3] ), .Y(n739) );
  NAND2X1 U1047 ( .A(n529), .B(\ab[7][3] ), .Y(n740) );
  NAND3X1 U1048 ( .A(n739), .B(n740), .C(n738), .Y(\CARRYB[7][3] ) );
  XOR2X1 U1049 ( .A(n528), .B(\ab[13][1] ), .Y(n837) );
  XOR2X1 U1050 ( .A(\SUMB[14][5] ), .B(n741), .Y(\SUMB[15][4] ) );
  NAND2X1 U1051 ( .A(\SUMB[14][5] ), .B(n270), .Y(n742) );
  NAND2X1 U1052 ( .A(\SUMB[14][5] ), .B(\ab[15][4] ), .Y(n743) );
  NAND2X1 U1053 ( .A(n270), .B(\ab[15][4] ), .Y(n744) );
  NAND3X1 U1054 ( .A(n744), .B(n742), .C(n743), .Y(\CARRYB[15][4] ) );
  XOR2X1 U1055 ( .A(n745), .B(\SUMB[11][8] ), .Y(\SUMB[12][7] ) );
  NAND2X1 U1056 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .Y(n746) );
  NAND2X1 U1057 ( .A(\ab[11][8] ), .B(\SUMB[10][9] ), .Y(n747) );
  NAND2X1 U1058 ( .A(\CARRYB[10][8] ), .B(\SUMB[10][9] ), .Y(n748) );
  NAND3X1 U1059 ( .A(n746), .B(n747), .C(n748), .Y(\CARRYB[11][8] ) );
  NAND2X1 U1060 ( .A(\ab[12][7] ), .B(n571), .Y(n749) );
  NAND2X1 U1061 ( .A(\SUMB[11][8] ), .B(\ab[12][7] ), .Y(n750) );
  NAND2X1 U1062 ( .A(n571), .B(\SUMB[11][8] ), .Y(n751) );
  NAND3X1 U1063 ( .A(n749), .B(n750), .C(n751), .Y(\CARRYB[12][7] ) );
  XOR2X1 U1064 ( .A(\ab[7][12] ), .B(n239), .Y(n752) );
  XOR2X1 U1065 ( .A(n752), .B(\SUMB[6][13] ), .Y(\SUMB[7][12] ) );
  XOR2X1 U1066 ( .A(\CARRYB[7][11] ), .B(\ab[8][11] ), .Y(n753) );
  XOR2X1 U1067 ( .A(n753), .B(\SUMB[7][12] ), .Y(\SUMB[8][11] ) );
  NAND2X1 U1068 ( .A(\ab[7][12] ), .B(n239), .Y(n754) );
  NAND2X1 U1069 ( .A(\ab[7][12] ), .B(\SUMB[6][13] ), .Y(n755) );
  NAND2X1 U1070 ( .A(n239), .B(\SUMB[6][13] ), .Y(n756) );
  NAND3X1 U1071 ( .A(n754), .B(n755), .C(n756), .Y(\CARRYB[7][12] ) );
  NAND2X1 U1072 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .Y(n757) );
  NAND2X1 U1073 ( .A(\ab[8][11] ), .B(\SUMB[7][12] ), .Y(n758) );
  NAND2X1 U1074 ( .A(\CARRYB[7][11] ), .B(\SUMB[7][12] ), .Y(n759) );
  NAND3X1 U1075 ( .A(n757), .B(n758), .C(n759), .Y(\CARRYB[8][11] ) );
  AND2X2 U1076 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Y(n760) );
  XOR2X1 U1077 ( .A(ZA), .B(n505), .Y(n761) );
  XOR2X1 U1078 ( .A(n607), .B(n761), .Y(\A1[13] ) );
  NAND2X1 U1079 ( .A(\SUMB[15][0] ), .B(ZA), .Y(n762) );
  NAND2X1 U1080 ( .A(\SUMB[15][0] ), .B(n505), .Y(n763) );
  NAND2X1 U1081 ( .A(ZA), .B(n505), .Y(n764) );
  NAND3X1 U1082 ( .A(n764), .B(n763), .C(n762), .Y(\A2[14] ) );
  NAND2X1 U1083 ( .A(\ab[11][3] ), .B(n159), .Y(n765) );
  NAND2X1 U1084 ( .A(\SUMB[10][4] ), .B(\ab[11][3] ), .Y(n766) );
  NAND2X1 U1085 ( .A(n159), .B(\SUMB[10][4] ), .Y(n767) );
  NAND3X1 U1086 ( .A(n765), .B(n766), .C(n767), .Y(\CARRYB[11][3] ) );
  NAND2X1 U1087 ( .A(n95), .B(\ab[12][2] ), .Y(n768) );
  NAND2X1 U1088 ( .A(\SUMB[11][3] ), .B(n95), .Y(n769) );
  NAND2X1 U1089 ( .A(\SUMB[11][3] ), .B(\ab[12][2] ), .Y(n770) );
  NAND3X1 U1090 ( .A(n768), .B(n770), .C(n769), .Y(\CARRYB[12][2] ) );
  XOR2X1 U1091 ( .A(\SUMB[4][8] ), .B(n771), .Y(\SUMB[5][7] ) );
  NAND2X1 U1092 ( .A(\ab[4][8] ), .B(n390), .Y(n772) );
  NAND2X1 U1093 ( .A(\SUMB[3][9] ), .B(\ab[4][8] ), .Y(n773) );
  NAND2X1 U1094 ( .A(n390), .B(\SUMB[3][9] ), .Y(n774) );
  NAND3X1 U1095 ( .A(n772), .B(n773), .C(n774), .Y(\CARRYB[4][8] ) );
  NAND2X1 U1096 ( .A(\ab[5][7] ), .B(n377), .Y(n775) );
  NAND2X1 U1097 ( .A(\SUMB[4][8] ), .B(\ab[5][7] ), .Y(n776) );
  NAND2X1 U1098 ( .A(\SUMB[4][8] ), .B(n377), .Y(n777) );
  NAND3X1 U1099 ( .A(n775), .B(n776), .C(n777), .Y(\CARRYB[5][7] ) );
  INVX1 U1100 ( .A(n1007), .Y(n1041) );
  NAND2X1 U1101 ( .A(\ab[9][7] ), .B(n467), .Y(n778) );
  NAND2X1 U1102 ( .A(\SUMB[8][8] ), .B(\ab[9][7] ), .Y(n779) );
  NAND2X1 U1103 ( .A(n467), .B(\SUMB[8][8] ), .Y(n780) );
  NAND3X1 U1104 ( .A(n778), .B(n779), .C(n780), .Y(\CARRYB[9][7] ) );
  NAND2X1 U1105 ( .A(n391), .B(\ab[10][6] ), .Y(n781) );
  NAND2X1 U1106 ( .A(\SUMB[9][7] ), .B(n391), .Y(n782) );
  NAND2X1 U1107 ( .A(\SUMB[9][7] ), .B(\ab[10][6] ), .Y(n783) );
  NAND3X1 U1108 ( .A(n781), .B(n782), .C(n783), .Y(\CARRYB[10][6] ) );
  INVX1 U1109 ( .A(n1011), .Y(n1039) );
  NAND2X1 U1110 ( .A(\ab[3][7] ), .B(n396), .Y(n784) );
  NAND2X1 U1111 ( .A(\SUMB[2][8] ), .B(\ab[3][7] ), .Y(n785) );
  NAND2X1 U1112 ( .A(\SUMB[2][8] ), .B(n396), .Y(n786) );
  NAND3X1 U1113 ( .A(n784), .B(n785), .C(n786), .Y(\CARRYB[3][7] ) );
  NAND2X1 U1114 ( .A(n446), .B(\ab[4][6] ), .Y(n787) );
  NAND2X1 U1115 ( .A(\SUMB[3][7] ), .B(\ab[4][6] ), .Y(n788) );
  NAND2X1 U1116 ( .A(\SUMB[3][7] ), .B(n446), .Y(n789) );
  NAND3X1 U1117 ( .A(n787), .B(n789), .C(n788), .Y(\CARRYB[4][6] ) );
  NAND2X1 U1118 ( .A(\SUMB[1][9] ), .B(n415), .Y(n790) );
  NAND2X1 U1119 ( .A(\ab[2][8] ), .B(n415), .Y(n791) );
  NAND2X1 U1120 ( .A(\SUMB[1][9] ), .B(\ab[2][8] ), .Y(n792) );
  NAND2X1 U1121 ( .A(\ab[10][5] ), .B(n93), .Y(n793) );
  NAND2X1 U1122 ( .A(\SUMB[9][6] ), .B(\ab[10][5] ), .Y(n794) );
  NAND2X1 U1123 ( .A(\SUMB[9][6] ), .B(n93), .Y(n795) );
  NAND3X1 U1124 ( .A(n794), .B(n793), .C(n795), .Y(\CARRYB[10][5] ) );
  NAND2X1 U1125 ( .A(\ab[11][4] ), .B(n971), .Y(n796) );
  NAND2X1 U1126 ( .A(\SUMB[10][5] ), .B(\ab[11][4] ), .Y(n797) );
  NAND2X1 U1127 ( .A(\SUMB[10][5] ), .B(n971), .Y(n798) );
  NAND3X1 U1128 ( .A(n796), .B(n797), .C(n798), .Y(\CARRYB[11][4] ) );
  NAND2X1 U1129 ( .A(\SUMB[8][7] ), .B(\CARRYB[8][6] ), .Y(n799) );
  NAND2X1 U1130 ( .A(\SUMB[8][7] ), .B(\ab[9][6] ), .Y(n800) );
  NAND2X1 U1131 ( .A(n45), .B(\ab[9][6] ), .Y(n801) );
  NAND3X1 U1132 ( .A(n801), .B(n799), .C(n800), .Y(\CARRYB[9][6] ) );
  AND2X2 U1133 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Y(n802) );
  XOR2X1 U1134 ( .A(n981), .B(n804), .Y(n883) );
  NAND2X1 U1135 ( .A(\ab[9][8] ), .B(n236), .Y(n805) );
  NAND2X1 U1136 ( .A(\SUMB[8][9] ), .B(\ab[9][8] ), .Y(n806) );
  NAND2X1 U1137 ( .A(n236), .B(\SUMB[8][9] ), .Y(n807) );
  NAND3X1 U1138 ( .A(n805), .B(n806), .C(n807), .Y(\CARRYB[9][8] ) );
  NAND2X1 U1139 ( .A(\ab[10][7] ), .B(n272), .Y(n808) );
  NAND2X1 U1140 ( .A(\SUMB[9][8] ), .B(\ab[10][7] ), .Y(n809) );
  NAND2X1 U1141 ( .A(\SUMB[9][8] ), .B(n272), .Y(n810) );
  NAND3X1 U1142 ( .A(n808), .B(n809), .C(n810), .Y(\CARRYB[10][7] ) );
  NAND2X1 U1143 ( .A(\SUMB[12][5] ), .B(n703), .Y(n812) );
  NAND2X1 U1144 ( .A(\SUMB[12][5] ), .B(\ab[13][4] ), .Y(n813) );
  NAND2X1 U1145 ( .A(n703), .B(\ab[13][4] ), .Y(n814) );
  NAND3X1 U1146 ( .A(n813), .B(n812), .C(n814), .Y(\CARRYB[13][4] ) );
  NAND2X1 U1147 ( .A(\SUMB[7][9] ), .B(n480), .Y(n815) );
  NAND2X1 U1148 ( .A(\SUMB[7][9] ), .B(\ab[8][8] ), .Y(n816) );
  NAND2X1 U1149 ( .A(n480), .B(\ab[8][8] ), .Y(n817) );
  NAND3X1 U1150 ( .A(n816), .B(n815), .C(n817), .Y(\CARRYB[8][8] ) );
  NAND2X1 U1151 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .Y(n818) );
  NAND2X1 U1152 ( .A(\ab[4][10] ), .B(\SUMB[3][11] ), .Y(n819) );
  NAND2X1 U1153 ( .A(\CARRYB[3][10] ), .B(\SUMB[3][11] ), .Y(n820) );
  NAND2X1 U1154 ( .A(n77), .B(\ab[5][10] ), .Y(n821) );
  NAND2X1 U1155 ( .A(\ab[5][10] ), .B(n112), .Y(n822) );
  NAND2X1 U1156 ( .A(n77), .B(n112), .Y(n823) );
  NAND3X1 U1157 ( .A(n821), .B(n822), .C(n823), .Y(\CARRYB[5][10] ) );
  NAND2X1 U1158 ( .A(\ab[12][6] ), .B(n273), .Y(n824) );
  NAND2X1 U1159 ( .A(\SUMB[11][7] ), .B(\ab[12][6] ), .Y(n825) );
  NAND2X1 U1160 ( .A(\SUMB[11][7] ), .B(n273), .Y(n826) );
  NAND3X1 U1161 ( .A(n824), .B(n825), .C(n826), .Y(\CARRYB[12][6] ) );
  NAND2X1 U1162 ( .A(\ab[13][5] ), .B(n82), .Y(n827) );
  NAND2X1 U1163 ( .A(\SUMB[12][6] ), .B(\ab[13][5] ), .Y(n828) );
  NAND2X1 U1164 ( .A(\SUMB[12][6] ), .B(n82), .Y(n829) );
  XOR2X1 U1165 ( .A(n345), .B(\ab[6][11] ), .Y(n830) );
  XOR2X1 U1166 ( .A(n830), .B(\SUMB[5][12] ), .Y(\SUMB[6][11] ) );
  NAND2X1 U1167 ( .A(\SUMB[5][12] ), .B(n345), .Y(n831) );
  NAND2X1 U1168 ( .A(\SUMB[5][12] ), .B(\ab[6][11] ), .Y(n832) );
  NAND2X1 U1169 ( .A(n345), .B(\ab[6][11] ), .Y(n833) );
  NAND3X1 U1170 ( .A(n832), .B(n831), .C(n833), .Y(\CARRYB[6][11] ) );
  NAND2X1 U1171 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(n834) );
  NAND2X1 U1172 ( .A(\CARRYB[7][9] ), .B(\ab[8][9] ), .Y(n835) );
  NAND2X1 U1173 ( .A(\SUMB[7][10] ), .B(\ab[8][9] ), .Y(n836) );
  NAND3X1 U1174 ( .A(n835), .B(n834), .C(n836), .Y(\CARRYB[8][9] ) );
  INVX1 U1175 ( .A(n1015), .Y(n1037) );
  NAND2X1 U1176 ( .A(\CARRYB[12][1] ), .B(\SUMB[12][2] ), .Y(n838) );
  NAND2X1 U1177 ( .A(\SUMB[12][2] ), .B(\ab[13][1] ), .Y(n839) );
  NAND2X1 U1178 ( .A(\CARRYB[12][1] ), .B(\ab[13][1] ), .Y(n840) );
  NAND3X1 U1179 ( .A(n839), .B(n838), .C(n840), .Y(\CARRYB[13][1] ) );
  INVX2 U1180 ( .A(\CARRYB[3][6] ), .Y(n841) );
  NAND2X1 U1181 ( .A(\ab[12][4] ), .B(n369), .Y(n842) );
  NAND2X1 U1182 ( .A(\SUMB[11][5] ), .B(\ab[12][4] ), .Y(n843) );
  NAND2X1 U1183 ( .A(\SUMB[11][5] ), .B(n369), .Y(n844) );
  NAND3X1 U1184 ( .A(n842), .B(n843), .C(n844), .Y(\CARRYB[12][4] ) );
  NAND2X1 U1185 ( .A(\CARRYB[12][3] ), .B(\ab[13][3] ), .Y(n845) );
  NAND2X1 U1186 ( .A(\ab[13][3] ), .B(\SUMB[12][4] ), .Y(n846) );
  NAND2X1 U1187 ( .A(\SUMB[12][4] ), .B(\CARRYB[12][3] ), .Y(n847) );
  NAND2X1 U1188 ( .A(\SUMB[3][13] ), .B(n346), .Y(n848) );
  NAND2X1 U1189 ( .A(\SUMB[3][13] ), .B(\ab[4][12] ), .Y(n849) );
  NAND2X1 U1190 ( .A(n346), .B(\ab[4][12] ), .Y(n850) );
  NAND3X1 U1191 ( .A(n849), .B(n848), .C(n850), .Y(\CARRYB[4][12] ) );
  XOR2X1 U1192 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .Y(n851) );
  XOR2X1 U1193 ( .A(n851), .B(\SUMB[4][12] ), .Y(\SUMB[5][11] ) );
  XOR2X1 U1194 ( .A(n852), .B(n18), .Y(\SUMB[6][10] ) );
  NAND2X1 U1195 ( .A(\ab[5][11] ), .B(n249), .Y(n853) );
  NAND2X1 U1196 ( .A(\SUMB[4][12] ), .B(\ab[5][11] ), .Y(n854) );
  NAND2X1 U1197 ( .A(\SUMB[4][12] ), .B(n249), .Y(n855) );
  NAND2X1 U1198 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .Y(n856) );
  NAND2X1 U1199 ( .A(\ab[6][10] ), .B(\SUMB[5][11] ), .Y(n857) );
  NAND2X1 U1200 ( .A(\CARRYB[5][10] ), .B(\SUMB[5][11] ), .Y(n858) );
  NAND3X1 U1201 ( .A(n856), .B(n857), .C(n858), .Y(\CARRYB[6][10] ) );
  NAND2X1 U1202 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .Y(n859) );
  NAND2X1 U1203 ( .A(\SUMB[3][10] ), .B(\ab[4][9] ), .Y(n860) );
  NAND2X1 U1204 ( .A(\CARRYB[3][9] ), .B(\SUMB[3][10] ), .Y(n861) );
  NAND3X1 U1205 ( .A(n860), .B(n859), .C(n861), .Y(\CARRYB[4][9] ) );
  NAND2X1 U1206 ( .A(\ab[5][8] ), .B(n601), .Y(n862) );
  NAND2X1 U1207 ( .A(\SUMB[4][9] ), .B(\ab[5][8] ), .Y(n863) );
  NAND2X1 U1208 ( .A(\SUMB[4][9] ), .B(n601), .Y(n864) );
  NAND3X1 U1209 ( .A(n862), .B(n863), .C(n864), .Y(\CARRYB[5][8] ) );
  NAND2X1 U1210 ( .A(\ab[8][6] ), .B(n318), .Y(n865) );
  NAND2X1 U1211 ( .A(\SUMB[7][7] ), .B(\ab[8][6] ), .Y(n866) );
  NAND2X1 U1212 ( .A(\SUMB[7][7] ), .B(n318), .Y(n867) );
  NAND3X1 U1213 ( .A(n865), .B(n866), .C(n867), .Y(\CARRYB[8][6] ) );
  NAND2X1 U1214 ( .A(\ab[9][5] ), .B(n600), .Y(n868) );
  NAND2X1 U1215 ( .A(\ab[9][5] ), .B(\SUMB[8][6] ), .Y(n869) );
  NAND2X1 U1216 ( .A(n600), .B(\SUMB[8][6] ), .Y(n870) );
  NAND3X1 U1217 ( .A(n868), .B(n869), .C(n870), .Y(\CARRYB[9][5] ) );
  XOR2X1 U1218 ( .A(n386), .B(\ab[14][0] ), .Y(n871) );
  XOR2X1 U1219 ( .A(n704), .B(n871), .Y(\A1[12] ) );
  NAND2X1 U1220 ( .A(\SUMB[13][1] ), .B(\CARRYB[13][0] ), .Y(n872) );
  NAND2X1 U1221 ( .A(\SUMB[13][1] ), .B(\ab[14][0] ), .Y(n873) );
  NAND2X1 U1222 ( .A(\CARRYB[13][0] ), .B(\ab[14][0] ), .Y(n874) );
  NAND3X1 U1223 ( .A(n874), .B(n872), .C(n873), .Y(\CARRYB[14][0] ) );
  NAND2X1 U1224 ( .A(\SUMB[7][5] ), .B(n543), .Y(n877) );
  NAND2X1 U1225 ( .A(\SUMB[7][5] ), .B(\ab[8][4] ), .Y(n878) );
  NAND2X1 U1226 ( .A(n543), .B(\ab[8][4] ), .Y(n879) );
  NAND3X1 U1227 ( .A(n879), .B(n877), .C(n878), .Y(\CARRYB[8][4] ) );
  NAND2X1 U1228 ( .A(\SUMB[7][6] ), .B(n278), .Y(n880) );
  NAND2X1 U1229 ( .A(\SUMB[7][6] ), .B(\ab[8][5] ), .Y(n881) );
  NAND2X1 U1230 ( .A(n278), .B(\ab[8][5] ), .Y(n882) );
  NAND3X1 U1231 ( .A(n882), .B(n881), .C(n880), .Y(\CARRYB[8][5] ) );
  XOR2X1 U1232 ( .A(\ab[13][0] ), .B(n388), .Y(n884) );
  XOR2X1 U1233 ( .A(n884), .B(n548), .Y(\A1[11] ) );
  NAND2X1 U1234 ( .A(\ab[12][1] ), .B(n982), .Y(n885) );
  NAND2X1 U1235 ( .A(\SUMB[11][2] ), .B(\ab[12][1] ), .Y(n886) );
  NAND2X1 U1236 ( .A(n982), .B(\SUMB[11][2] ), .Y(n887) );
  NAND3X1 U1237 ( .A(n885), .B(n887), .C(n886), .Y(\CARRYB[12][1] ) );
  NAND2X1 U1238 ( .A(\CARRYB[12][0] ), .B(\ab[13][0] ), .Y(n888) );
  NAND2X1 U1239 ( .A(\ab[13][0] ), .B(\SUMB[12][1] ), .Y(n889) );
  NAND2X1 U1240 ( .A(\CARRYB[12][0] ), .B(\SUMB[12][1] ), .Y(n890) );
  NAND3X1 U1241 ( .A(n889), .B(n890), .C(n888), .Y(\CARRYB[13][0] ) );
  NAND2X1 U1242 ( .A(n538), .B(n301), .Y(n891) );
  NAND2X1 U1243 ( .A(\SUMB[2][9] ), .B(n538), .Y(n892) );
  NAND2X1 U1244 ( .A(\SUMB[2][9] ), .B(n301), .Y(n893) );
  NAND3X1 U1245 ( .A(n891), .B(n892), .C(n893), .Y(\CARRYB[3][8] ) );
  NAND2X1 U1246 ( .A(n475), .B(\ab[4][7] ), .Y(n894) );
  NAND2X1 U1247 ( .A(\ab[4][7] ), .B(\SUMB[3][8] ), .Y(n895) );
  NAND2X1 U1248 ( .A(\SUMB[3][8] ), .B(n475), .Y(n896) );
  NAND3X1 U1249 ( .A(n894), .B(n896), .C(n895), .Y(\CARRYB[4][7] ) );
  XOR2X1 U1250 ( .A(\SUMB[6][8] ), .B(n897), .Y(\SUMB[7][7] ) );
  NAND2X1 U1251 ( .A(\ab[6][8] ), .B(n393), .Y(n898) );
  NAND2X1 U1252 ( .A(\SUMB[5][9] ), .B(\ab[6][8] ), .Y(n899) );
  NAND2X1 U1253 ( .A(\SUMB[5][9] ), .B(n393), .Y(n900) );
  NAND3X1 U1254 ( .A(n898), .B(n899), .C(n900), .Y(\CARRYB[6][8] ) );
  NAND2X1 U1255 ( .A(n44), .B(\ab[7][7] ), .Y(n901) );
  NAND2X1 U1256 ( .A(\SUMB[6][8] ), .B(\ab[7][7] ), .Y(n902) );
  NAND2X1 U1257 ( .A(\SUMB[6][8] ), .B(n256), .Y(n903) );
  NAND3X1 U1258 ( .A(n901), .B(n902), .C(n903), .Y(\CARRYB[7][7] ) );
  INVX1 U1259 ( .A(n507), .Y(n1042) );
  AND2X2 U1260 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(n904) );
  INVX2 U1261 ( .A(n1002), .Y(n1003) );
  INVX2 U1262 ( .A(B[7]), .Y(n1002) );
  INVX1 U1263 ( .A(n905), .Y(n1043) );
  INVX4 U1264 ( .A(n1000), .Y(n969) );
  AND2X2 U1265 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(n906) );
  NAND2X1 U1266 ( .A(n655), .B(ZB), .Y(n907) );
  NAND2X1 U1267 ( .A(\ab[3][12] ), .B(n271), .Y(n908) );
  NAND2X1 U1268 ( .A(\SUMB[2][13] ), .B(\ab[3][12] ), .Y(n909) );
  NAND2X1 U1269 ( .A(n271), .B(\SUMB[2][13] ), .Y(n910) );
  NAND3X1 U1270 ( .A(n908), .B(n909), .C(n910), .Y(\CARRYB[3][12] ) );
  NAND2X1 U1271 ( .A(\ab[4][11] ), .B(n582), .Y(n911) );
  NAND2X1 U1272 ( .A(\SUMB[3][12] ), .B(\ab[4][11] ), .Y(n912) );
  NAND2X1 U1273 ( .A(\SUMB[3][12] ), .B(n582), .Y(n913) );
  NAND3X1 U1274 ( .A(n911), .B(n912), .C(n913), .Y(\CARRYB[4][11] ) );
  XOR2X1 U1275 ( .A(\SUMB[1][14] ), .B(n914), .Y(\SUMB[2][13] ) );
  NAND2X1 U1276 ( .A(\SUMB[1][14] ), .B(\ab[2][13] ), .Y(n915) );
  NAND2X1 U1277 ( .A(\SUMB[1][14] ), .B(n246), .Y(n916) );
  NAND2X1 U1278 ( .A(\ab[2][13] ), .B(n246), .Y(n917) );
  NAND3X1 U1279 ( .A(n916), .B(n915), .C(n917), .Y(\CARRYB[2][13] ) );
  XOR2X1 U1280 ( .A(n918), .B(n76), .Y(\SUMB[14][1] ) );
  NAND2X1 U1281 ( .A(\ab[13][2] ), .B(n398), .Y(n919) );
  NAND2X1 U1282 ( .A(\SUMB[12][3] ), .B(\ab[13][2] ), .Y(n920) );
  NAND2X1 U1283 ( .A(\SUMB[12][3] ), .B(n398), .Y(n921) );
  NAND3X1 U1284 ( .A(n919), .B(n921), .C(n920), .Y(\CARRYB[13][2] ) );
  NAND2X1 U1285 ( .A(\ab[14][1] ), .B(n87), .Y(n922) );
  NAND2X1 U1286 ( .A(\SUMB[13][2] ), .B(\ab[14][1] ), .Y(n923) );
  NAND2X1 U1287 ( .A(\SUMB[13][2] ), .B(n87), .Y(n924) );
  NAND3X1 U1288 ( .A(n922), .B(n923), .C(n924), .Y(\CARRYB[14][1] ) );
  NAND2X1 U1289 ( .A(\ab[6][5] ), .B(n663), .Y(n925) );
  NAND2X1 U1290 ( .A(\SUMB[5][6] ), .B(\ab[6][5] ), .Y(n926) );
  NAND2X1 U1291 ( .A(\SUMB[5][6] ), .B(n663), .Y(n927) );
  NAND3X1 U1292 ( .A(n926), .B(n925), .C(n927), .Y(\CARRYB[6][5] ) );
  NAND2X1 U1293 ( .A(n14), .B(\ab[7][4] ), .Y(n928) );
  NAND2X1 U1294 ( .A(\SUMB[6][5] ), .B(\ab[7][4] ), .Y(n929) );
  NAND2X1 U1295 ( .A(n14), .B(\SUMB[6][5] ), .Y(n930) );
  NAND3X1 U1296 ( .A(n928), .B(n929), .C(n930), .Y(\CARRYB[7][4] ) );
  NAND2X1 U1297 ( .A(\SUMB[9][3] ), .B(n15), .Y(n931) );
  NAND2X1 U1298 ( .A(\SUMB[9][3] ), .B(\ab[10][2] ), .Y(n932) );
  NAND2X1 U1299 ( .A(n15), .B(\ab[10][2] ), .Y(n933) );
  NAND3X1 U1300 ( .A(n932), .B(n931), .C(n933), .Y(\CARRYB[10][2] ) );
  XOR2X1 U1301 ( .A(\ab[5][2] ), .B(n164), .Y(n935) );
  XOR2X1 U1302 ( .A(n935), .B(n321), .Y(\SUMB[5][2] ) );
  NAND2X1 U1303 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .Y(n936) );
  NAND2X1 U1304 ( .A(\ab[4][3] ), .B(\SUMB[3][4] ), .Y(n937) );
  NAND2X1 U1305 ( .A(\CARRYB[3][3] ), .B(\SUMB[3][4] ), .Y(n938) );
  NAND3X1 U1306 ( .A(n936), .B(n937), .C(n938), .Y(\CARRYB[4][3] ) );
  NAND2X1 U1307 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .Y(n939) );
  NAND2X1 U1308 ( .A(\ab[5][2] ), .B(\SUMB[4][3] ), .Y(n940) );
  NAND2X1 U1309 ( .A(\CARRYB[4][2] ), .B(\SUMB[4][3] ), .Y(n941) );
  NAND3X1 U1310 ( .A(n939), .B(n940), .C(n941), .Y(\CARRYB[5][2] ) );
  NAND2X1 U1311 ( .A(\ab[2][4] ), .B(n654), .Y(n942) );
  NAND2X1 U1312 ( .A(\ab[2][4] ), .B(\SUMB[1][5] ), .Y(n943) );
  NAND2X1 U1313 ( .A(n654), .B(\SUMB[1][5] ), .Y(n944) );
  NAND3X1 U1314 ( .A(n942), .B(n943), .C(n944), .Y(\CARRYB[2][4] ) );
  NAND2X1 U1315 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .Y(n945) );
  NAND2X1 U1316 ( .A(\ab[3][3] ), .B(\SUMB[2][4] ), .Y(n946) );
  NAND2X1 U1317 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n947) );
  NAND3X1 U1318 ( .A(n945), .B(n946), .C(n947), .Y(\CARRYB[3][3] ) );
  XOR2X1 U1319 ( .A(n457), .B(\ab[6][3] ), .Y(n948) );
  XOR2X1 U1320 ( .A(n526), .B(n948), .Y(\SUMB[6][3] ) );
  NAND2X1 U1321 ( .A(\SUMB[5][4] ), .B(\CARRYB[5][3] ), .Y(n949) );
  NAND2X1 U1322 ( .A(\SUMB[5][4] ), .B(\ab[6][3] ), .Y(n950) );
  NAND2X1 U1323 ( .A(\CARRYB[5][3] ), .B(\ab[6][3] ), .Y(n951) );
  NAND3X1 U1324 ( .A(n950), .B(n949), .C(n951), .Y(\CARRYB[6][3] ) );
  INVX2 U1325 ( .A(n999), .Y(n973) );
  BUFX4 U1326 ( .A(\CARRYB[2][0] ), .Y(n968) );
  AND2X2 U1327 ( .A(\SUMB[15][2] ), .B(\CARRYB[15][1] ), .Y(n953) );
  AND2X2 U1328 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n958) );
  AND2X2 U1329 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n959) );
  AND2X2 U1330 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n960) );
  NOR2X1 U1331 ( .A(n999), .B(n655), .Y(n962) );
  INVX2 U1332 ( .A(A[13]), .Y(n1054) );
  INVX2 U1333 ( .A(ZA), .Y(n1052) );
  INVX2 U1334 ( .A(A[14]), .Y(n1053) );
  INVX2 U1335 ( .A(A[4]), .Y(n1023) );
  INVX2 U1336 ( .A(A[5]), .Y(n1025) );
  INVX2 U1337 ( .A(A[6]), .Y(n1027) );
  INVX2 U1338 ( .A(A[7]), .Y(n1029) );
  INVX2 U1339 ( .A(A[8]), .Y(n1031) );
  INVX2 U1340 ( .A(A[9]), .Y(n1033) );
  INVX2 U1341 ( .A(A[10]), .Y(n1035) );
  XOR2X1 U1342 ( .A(\CARRYB[15][0] ), .B(\SUMB[15][1] ), .Y(\A1[14] ) );
  XOR2X1 U1343 ( .A(\SUMB[15][2] ), .B(\CARRYB[15][1] ), .Y(\A1[15] ) );
  XOR2X1 U1344 ( .A(\SUMB[15][4] ), .B(\CARRYB[15][3] ), .Y(\A1[17] ) );
  XOR2X1 U1345 ( .A(\SUMB[15][6] ), .B(\CARRYB[15][5] ), .Y(\A1[19] ) );
  NAND2X1 U1346 ( .A(\SUMB[15][7] ), .B(\CARRYB[15][6] ), .Y(n963) );
  INVX2 U1347 ( .A(n963), .Y(\A2[21] ) );
  XOR2X1 U1348 ( .A(\SUMB[15][8] ), .B(\CARRYB[15][7] ), .Y(\A1[21] ) );
  NAND2X1 U1349 ( .A(\SUMB[15][8] ), .B(\CARRYB[15][7] ), .Y(n964) );
  INVX2 U1350 ( .A(n964), .Y(\A2[22] ) );
  XOR2X1 U1351 ( .A(\SUMB[15][9] ), .B(\CARRYB[15][8] ), .Y(\A1[22] ) );
  XOR2X1 U1352 ( .A(\SUMB[15][10] ), .B(\CARRYB[15][9] ), .Y(\A1[23] ) );
  XOR2X1 U1353 ( .A(\SUMB[15][11] ), .B(\CARRYB[15][10] ), .Y(\A1[24] ) );
  XOR2X1 U1354 ( .A(\SUMB[15][12] ), .B(\CARRYB[15][11] ), .Y(\A1[25] ) );
  XOR2X1 U1355 ( .A(\SUMB[15][13] ), .B(\CARRYB[15][12] ), .Y(\A1[26] ) );
  XOR2X1 U1356 ( .A(\SUMB[15][14] ), .B(\CARRYB[15][13] ), .Y(\A1[27] ) );
  XOR2X1 U1357 ( .A(\SUMB[15][15] ), .B(\CARRYB[15][14] ), .Y(\A1[28] ) );
  XOR2X1 U1358 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U1359 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  NAND2X1 U1360 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n965) );
  INVX2 U1361 ( .A(n965), .Y(\CARRYB[1][1] ) );
  XOR2X1 U1362 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U1363 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U1364 ( .A(n962), .B(\ab[1][4] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U1365 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U1366 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U1367 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(\SUMB[1][7] ) );
  XOR2X1 U1368 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(\SUMB[1][8] ) );
  XOR2X1 U1369 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(\SUMB[1][11] ) );
  XOR2X1 U1370 ( .A(n96), .B(\ab[1][12] ), .Y(\SUMB[1][12] ) );
  NAND2X1 U1371 ( .A(\ab[0][14] ), .B(n139), .Y(n966) );
  XOR2X1 U1372 ( .A(\ab[1][14] ), .B(n984), .Y(\SUMB[1][14] ) );
  BUFX4 U1373 ( .A(\CARRYB[10][0] ), .Y(n967) );
  INVX2 U1374 ( .A(n1000), .Y(n1001) );
  INVX2 U1375 ( .A(B[6]), .Y(n1000) );
  INVX1 U1376 ( .A(n969), .Y(n1044) );
  INVX2 U1377 ( .A(\CARRYB[10][4] ), .Y(n970) );
  INVX1 U1378 ( .A(n999), .Y(n972) );
  INVX2 U1379 ( .A(B[5]), .Y(n999) );
  INVX2 U1380 ( .A(n989), .Y(n990) );
  INVX1 U1381 ( .A(n973), .Y(n1045) );
  INVX2 U1382 ( .A(\CARRYB[2][4] ), .Y(n975) );
  INVX2 U1383 ( .A(n993), .Y(n976) );
  INVX2 U1384 ( .A(n993), .Y(n994) );
  INVX2 U1385 ( .A(B[2]), .Y(n993) );
  INVX2 U1386 ( .A(n997), .Y(n998) );
  INVX2 U1387 ( .A(n995), .Y(n978) );
  INVX2 U1388 ( .A(n995), .Y(n996) );
  INVX2 U1389 ( .A(B[3]), .Y(n995) );
  INVX1 U1390 ( .A(n977), .Y(n1046) );
  INVX1 U1391 ( .A(n978), .Y(n1047) );
  INVX2 U1392 ( .A(n991), .Y(n992) );
  INVX2 U1393 ( .A(B[1]), .Y(n991) );
  INVX1 U1394 ( .A(n976), .Y(n1048) );
  INVX1 U1395 ( .A(n980), .Y(n1049) );
  INVX2 U1396 ( .A(n1016), .Y(n985) );
  INVX2 U1397 ( .A(\CARRYB[11][1] ), .Y(n981) );
  INVX2 U1398 ( .A(\CARRYB[2][3] ), .Y(n983) );
  INVX4 U1399 ( .A(A[1]), .Y(n1017) );
  INVX2 U1400 ( .A(\CARRYB[2][2] ), .Y(n986) );
  INVX8 U1401 ( .A(n1014), .Y(n1015) );
  INVX8 U1402 ( .A(n1021), .Y(n1022) );
  INVX8 U1403 ( .A(n1023), .Y(n1024) );
  INVX8 U1404 ( .A(n1025), .Y(n1026) );
  INVX8 U1405 ( .A(n1027), .Y(n1028) );
  INVX8 U1406 ( .A(n1029), .Y(n1030) );
  INVX8 U1407 ( .A(n1031), .Y(n1032) );
  INVX8 U1408 ( .A(n1033), .Y(n1034) );
  INVX8 U1409 ( .A(n1035), .Y(n1036) );
  AND2X2 U1410 ( .A(n1018), .B(B[14]), .Y(\ab[1][14] ) );
  AND2X2 U1411 ( .A(B[14]), .B(n401), .Y(\ab[0][14] ) );
  AND2X2 U1412 ( .A(n1018), .B(B[12]), .Y(\ab[1][12] ) );
  AND2X2 U1413 ( .A(B[12]), .B(n531), .Y(\ab[0][12] ) );
  AND2X2 U1414 ( .A(n423), .B(B[10]), .Y(\ab[1][10] ) );
  AND2X2 U1415 ( .A(n531), .B(B[10]), .Y(\ab[0][10] ) );
  AND2X2 U1416 ( .A(B[9]), .B(n531), .Y(\ab[0][9] ) );
  AND2X2 U1417 ( .A(n1018), .B(B[8]), .Y(\ab[1][8] ) );
  AND2X2 U1418 ( .A(n985), .B(B[8]), .Y(\ab[0][8] ) );
  AND2X2 U1419 ( .A(n1003), .B(n423), .Y(\ab[1][7] ) );
  AND2X2 U1420 ( .A(n1003), .B(n985), .Y(\ab[0][7] ) );
  AND2X2 U1421 ( .A(n1018), .B(n1001), .Y(\ab[1][6] ) );
  AND2X2 U1422 ( .A(n1001), .B(n402), .Y(\ab[0][6] ) );
  AND2X2 U1423 ( .A(B[5]), .B(n1018), .Y(\ab[1][5] ) );
  AND2X2 U1424 ( .A(n1018), .B(n998), .Y(\ab[1][4] ) );
  AND2X2 U1425 ( .A(n998), .B(n402), .Y(\ab[0][4] ) );
  AND2X2 U1426 ( .A(n1018), .B(n996), .Y(\ab[1][3] ) );
  AND2X2 U1427 ( .A(n996), .B(n401), .Y(\ab[0][3] ) );
  AND2X2 U1428 ( .A(n994), .B(n9), .Y(\ab[1][2] ) );
  AND2X2 U1429 ( .A(n994), .B(n402), .Y(\ab[0][2] ) );
  AND2X2 U1430 ( .A(n1018), .B(n992), .Y(\ab[1][1] ) );
  AND2X2 U1431 ( .A(n992), .B(n402), .Y(\ab[0][1] ) );
  AND2X2 U1432 ( .A(n9), .B(n990), .Y(\ab[1][0] ) );
  NOR2X1 U1433 ( .A(n1018), .B(n1051), .Y(\ab[1][15] ) );
  AND2X2 U1434 ( .A(n4), .B(n1013), .Y(\ab[2][13] ) );
  AND2X2 U1435 ( .A(n5), .B(n1011), .Y(\ab[2][12] ) );
  AND2X2 U1436 ( .A(n5), .B(n1009), .Y(\ab[2][11] ) );
  AND2X2 U1437 ( .A(n1020), .B(n1007), .Y(\ab[2][10] ) );
  AND2X2 U1438 ( .A(n1020), .B(B[9]), .Y(\ab[2][9] ) );
  AND2X2 U1439 ( .A(n1020), .B(B[8]), .Y(\ab[2][8] ) );
  AND2X2 U1440 ( .A(n4), .B(n969), .Y(\ab[2][6] ) );
  AND2X2 U1441 ( .A(n5), .B(n973), .Y(\ab[2][5] ) );
  AND2X2 U1442 ( .A(n4), .B(n977), .Y(\ab[2][4] ) );
  AND2X2 U1443 ( .A(n10), .B(n978), .Y(\ab[2][3] ) );
  AND2X2 U1444 ( .A(n10), .B(n976), .Y(\ab[2][2] ) );
  AND2X2 U1445 ( .A(n5), .B(n980), .Y(\ab[2][1] ) );
  AND2X2 U1446 ( .A(n5), .B(n974), .Y(\ab[2][0] ) );
  AND2X2 U1447 ( .A(n1022), .B(n1015), .Y(\ab[3][14] ) );
  NOR2X1 U1448 ( .A(n4), .B(n1051), .Y(\ab[2][15] ) );
  AND2X2 U1449 ( .A(n1022), .B(n1013), .Y(\ab[3][13] ) );
  AND2X2 U1450 ( .A(n1022), .B(n1011), .Y(\ab[3][12] ) );
  AND2X2 U1451 ( .A(n1022), .B(n1009), .Y(\ab[3][11] ) );
  AND2X2 U1452 ( .A(n1022), .B(n1007), .Y(\ab[3][10] ) );
  AND2X2 U1453 ( .A(n1022), .B(n507), .Y(\ab[3][9] ) );
  AND2X2 U1454 ( .A(n1022), .B(n905), .Y(\ab[3][7] ) );
  AND2X2 U1455 ( .A(n1022), .B(n969), .Y(\ab[3][6] ) );
  AND2X2 U1456 ( .A(n1022), .B(n972), .Y(\ab[3][5] ) );
  AND2X2 U1457 ( .A(n1022), .B(n977), .Y(\ab[3][4] ) );
  AND2X2 U1458 ( .A(n1022), .B(n978), .Y(\ab[3][3] ) );
  AND2X2 U1459 ( .A(n1022), .B(n976), .Y(\ab[3][2] ) );
  AND2X2 U1460 ( .A(n1022), .B(n980), .Y(\ab[3][1] ) );
  AND2X2 U1461 ( .A(n1022), .B(n974), .Y(\ab[3][0] ) );
  AND2X2 U1462 ( .A(n1024), .B(n1015), .Y(\ab[4][14] ) );
  NOR2X1 U1463 ( .A(n1022), .B(n1051), .Y(\ab[3][15] ) );
  AND2X2 U1464 ( .A(n1024), .B(n1013), .Y(\ab[4][13] ) );
  AND2X2 U1465 ( .A(n1024), .B(n1011), .Y(\ab[4][12] ) );
  AND2X2 U1466 ( .A(n1024), .B(n1009), .Y(\ab[4][11] ) );
  AND2X2 U1467 ( .A(n1024), .B(n1007), .Y(\ab[4][10] ) );
  AND2X2 U1468 ( .A(n1024), .B(n507), .Y(\ab[4][9] ) );
  AND2X2 U1469 ( .A(n1024), .B(n1005), .Y(\ab[4][8] ) );
  AND2X2 U1470 ( .A(n1024), .B(n905), .Y(\ab[4][7] ) );
  AND2X2 U1471 ( .A(n1024), .B(n969), .Y(\ab[4][6] ) );
  AND2X2 U1472 ( .A(n1024), .B(n973), .Y(\ab[4][5] ) );
  AND2X2 U1473 ( .A(n1024), .B(n977), .Y(\ab[4][4] ) );
  AND2X2 U1474 ( .A(n1024), .B(n978), .Y(\ab[4][3] ) );
  AND2X2 U1475 ( .A(n1024), .B(n976), .Y(\ab[4][2] ) );
  AND2X2 U1476 ( .A(n1024), .B(n980), .Y(\ab[4][1] ) );
  AND2X2 U1477 ( .A(n1024), .B(n974), .Y(\ab[4][0] ) );
  AND2X2 U1478 ( .A(n1026), .B(n1015), .Y(\ab[5][14] ) );
  NOR2X1 U1479 ( .A(n1024), .B(n1051), .Y(\ab[4][15] ) );
  AND2X2 U1480 ( .A(n1026), .B(n1013), .Y(\ab[5][13] ) );
  AND2X2 U1481 ( .A(n1026), .B(n1011), .Y(\ab[5][12] ) );
  AND2X2 U1482 ( .A(n1026), .B(n163), .Y(\ab[5][11] ) );
  AND2X2 U1483 ( .A(n1026), .B(n1007), .Y(\ab[5][10] ) );
  AND2X2 U1484 ( .A(n1026), .B(n507), .Y(\ab[5][9] ) );
  AND2X2 U1485 ( .A(n1026), .B(n1005), .Y(\ab[5][8] ) );
  AND2X2 U1486 ( .A(n1026), .B(n905), .Y(\ab[5][7] ) );
  AND2X2 U1487 ( .A(n1026), .B(n969), .Y(\ab[5][6] ) );
  AND2X2 U1488 ( .A(n1026), .B(n972), .Y(\ab[5][5] ) );
  AND2X2 U1489 ( .A(n1026), .B(n977), .Y(\ab[5][4] ) );
  AND2X2 U1490 ( .A(n1026), .B(n978), .Y(\ab[5][3] ) );
  AND2X2 U1491 ( .A(n1026), .B(n976), .Y(\ab[5][2] ) );
  AND2X2 U1492 ( .A(n1026), .B(n980), .Y(\ab[5][1] ) );
  AND2X2 U1493 ( .A(n1026), .B(n974), .Y(\ab[5][0] ) );
  AND2X2 U1494 ( .A(n1028), .B(n1015), .Y(\ab[6][14] ) );
  NOR2X1 U1495 ( .A(n1026), .B(n1051), .Y(\ab[5][15] ) );
  AND2X2 U1496 ( .A(n1028), .B(n1013), .Y(\ab[6][13] ) );
  AND2X2 U1497 ( .A(n1028), .B(n1011), .Y(\ab[6][12] ) );
  AND2X2 U1498 ( .A(n1028), .B(n163), .Y(\ab[6][11] ) );
  AND2X2 U1499 ( .A(n1028), .B(n1007), .Y(\ab[6][10] ) );
  AND2X2 U1500 ( .A(n1028), .B(n507), .Y(\ab[6][9] ) );
  AND2X2 U1501 ( .A(n1028), .B(n1005), .Y(\ab[6][8] ) );
  AND2X2 U1502 ( .A(n1028), .B(n905), .Y(\ab[6][7] ) );
  AND2X2 U1503 ( .A(n1028), .B(n969), .Y(\ab[6][6] ) );
  AND2X2 U1504 ( .A(n1028), .B(n973), .Y(\ab[6][5] ) );
  AND2X2 U1505 ( .A(n1028), .B(n977), .Y(\ab[6][4] ) );
  AND2X2 U1506 ( .A(n1028), .B(n978), .Y(\ab[6][3] ) );
  AND2X2 U1507 ( .A(n1028), .B(n976), .Y(\ab[6][2] ) );
  AND2X2 U1508 ( .A(n1028), .B(n980), .Y(\ab[6][1] ) );
  AND2X2 U1509 ( .A(n1028), .B(n974), .Y(\ab[6][0] ) );
  AND2X2 U1510 ( .A(n1030), .B(n1015), .Y(\ab[7][14] ) );
  NOR2X1 U1511 ( .A(n1028), .B(n1051), .Y(\ab[6][15] ) );
  AND2X2 U1512 ( .A(n1030), .B(n1013), .Y(\ab[7][13] ) );
  AND2X2 U1513 ( .A(n1030), .B(n1011), .Y(\ab[7][12] ) );
  AND2X2 U1514 ( .A(n1030), .B(n163), .Y(\ab[7][11] ) );
  AND2X2 U1515 ( .A(n1030), .B(n1007), .Y(\ab[7][10] ) );
  AND2X2 U1516 ( .A(n1030), .B(n507), .Y(\ab[7][9] ) );
  AND2X2 U1517 ( .A(n1030), .B(n1005), .Y(\ab[7][8] ) );
  AND2X2 U1518 ( .A(n1030), .B(n905), .Y(\ab[7][7] ) );
  AND2X2 U1519 ( .A(n1030), .B(n969), .Y(\ab[7][6] ) );
  AND2X2 U1520 ( .A(n1030), .B(n972), .Y(\ab[7][5] ) );
  AND2X2 U1521 ( .A(n1030), .B(n977), .Y(\ab[7][4] ) );
  AND2X2 U1522 ( .A(n1030), .B(n978), .Y(\ab[7][3] ) );
  AND2X2 U1523 ( .A(n1030), .B(n976), .Y(\ab[7][2] ) );
  AND2X2 U1524 ( .A(n1030), .B(n980), .Y(\ab[7][1] ) );
  AND2X2 U1525 ( .A(n1030), .B(n974), .Y(\ab[7][0] ) );
  AND2X2 U1526 ( .A(n1032), .B(n1015), .Y(\ab[8][14] ) );
  NOR2X1 U1527 ( .A(n1030), .B(n1051), .Y(\ab[7][15] ) );
  AND2X2 U1528 ( .A(n1032), .B(n1013), .Y(\ab[8][13] ) );
  AND2X2 U1529 ( .A(n1032), .B(n1011), .Y(\ab[8][12] ) );
  AND2X2 U1530 ( .A(n1032), .B(n163), .Y(\ab[8][11] ) );
  AND2X2 U1531 ( .A(n1032), .B(n1007), .Y(\ab[8][10] ) );
  AND2X2 U1532 ( .A(n1032), .B(n507), .Y(\ab[8][9] ) );
  AND2X2 U1533 ( .A(n1032), .B(n1005), .Y(\ab[8][8] ) );
  AND2X2 U1534 ( .A(n1032), .B(n905), .Y(\ab[8][7] ) );
  AND2X2 U1535 ( .A(n1032), .B(n969), .Y(\ab[8][6] ) );
  AND2X2 U1536 ( .A(n1032), .B(n973), .Y(\ab[8][5] ) );
  AND2X2 U1537 ( .A(n1032), .B(n977), .Y(\ab[8][4] ) );
  AND2X2 U1538 ( .A(n1032), .B(n978), .Y(\ab[8][3] ) );
  AND2X2 U1539 ( .A(n1032), .B(n976), .Y(\ab[8][2] ) );
  AND2X2 U1540 ( .A(n1032), .B(n980), .Y(\ab[8][1] ) );
  AND2X2 U1541 ( .A(n1032), .B(n974), .Y(\ab[8][0] ) );
  AND2X2 U1542 ( .A(n1034), .B(n1015), .Y(\ab[9][14] ) );
  NOR2X1 U1543 ( .A(n1032), .B(n1051), .Y(\ab[8][15] ) );
  AND2X2 U1544 ( .A(n1034), .B(n1013), .Y(\ab[9][13] ) );
  AND2X2 U1545 ( .A(n1034), .B(n1011), .Y(\ab[9][12] ) );
  AND2X2 U1546 ( .A(n1034), .B(n163), .Y(\ab[9][11] ) );
  AND2X2 U1547 ( .A(n1034), .B(n1007), .Y(\ab[9][10] ) );
  AND2X2 U1548 ( .A(n1034), .B(n507), .Y(\ab[9][9] ) );
  AND2X2 U1549 ( .A(n1034), .B(n1005), .Y(\ab[9][8] ) );
  AND2X2 U1550 ( .A(n1034), .B(n905), .Y(\ab[9][7] ) );
  AND2X2 U1551 ( .A(n1034), .B(n969), .Y(\ab[9][6] ) );
  AND2X2 U1552 ( .A(n1034), .B(n972), .Y(\ab[9][5] ) );
  AND2X2 U1553 ( .A(n1034), .B(n977), .Y(\ab[9][4] ) );
  AND2X2 U1554 ( .A(n1034), .B(n978), .Y(\ab[9][3] ) );
  AND2X2 U1555 ( .A(n1034), .B(n976), .Y(\ab[9][2] ) );
  AND2X2 U1556 ( .A(n1034), .B(n980), .Y(\ab[9][1] ) );
  AND2X2 U1557 ( .A(n1034), .B(n974), .Y(\ab[9][0] ) );
  AND2X2 U1558 ( .A(n1036), .B(n1015), .Y(\ab[10][14] ) );
  NOR2X1 U1559 ( .A(n1034), .B(n1051), .Y(\ab[9][15] ) );
  AND2X2 U1560 ( .A(n1036), .B(n1013), .Y(\ab[10][13] ) );
  AND2X2 U1561 ( .A(n1036), .B(n1011), .Y(\ab[10][12] ) );
  AND2X2 U1562 ( .A(n1036), .B(n163), .Y(\ab[10][11] ) );
  AND2X2 U1563 ( .A(n1036), .B(n1007), .Y(\ab[10][10] ) );
  AND2X2 U1564 ( .A(n1036), .B(n507), .Y(\ab[10][9] ) );
  AND2X2 U1565 ( .A(n1036), .B(n1005), .Y(\ab[10][8] ) );
  AND2X2 U1566 ( .A(n1036), .B(n905), .Y(\ab[10][7] ) );
  AND2X2 U1567 ( .A(n1036), .B(n969), .Y(\ab[10][6] ) );
  AND2X2 U1568 ( .A(n1036), .B(n973), .Y(\ab[10][5] ) );
  AND2X2 U1569 ( .A(n1036), .B(n977), .Y(\ab[10][4] ) );
  AND2X2 U1570 ( .A(n1036), .B(n978), .Y(\ab[10][3] ) );
  AND2X2 U1571 ( .A(n1036), .B(n976), .Y(\ab[10][2] ) );
  AND2X2 U1572 ( .A(n1036), .B(n980), .Y(\ab[10][1] ) );
  AND2X2 U1573 ( .A(n1036), .B(n974), .Y(\ab[10][0] ) );
  AND2X2 U1574 ( .A(A[11]), .B(n1015), .Y(\ab[11][14] ) );
  NOR2X1 U1575 ( .A(n1036), .B(n1051), .Y(\ab[10][15] ) );
  AND2X2 U1576 ( .A(A[11]), .B(n1013), .Y(\ab[11][13] ) );
  AND2X2 U1577 ( .A(A[11]), .B(n1011), .Y(\ab[11][12] ) );
  AND2X2 U1578 ( .A(A[11]), .B(n163), .Y(\ab[11][11] ) );
  AND2X2 U1579 ( .A(A[11]), .B(n1007), .Y(\ab[11][10] ) );
  AND2X2 U1580 ( .A(A[11]), .B(n507), .Y(\ab[11][9] ) );
  AND2X2 U1581 ( .A(A[11]), .B(n1005), .Y(\ab[11][8] ) );
  AND2X2 U1582 ( .A(A[11]), .B(n905), .Y(\ab[11][7] ) );
  AND2X2 U1583 ( .A(A[11]), .B(n969), .Y(\ab[11][6] ) );
  AND2X2 U1584 ( .A(A[11]), .B(n972), .Y(\ab[11][5] ) );
  AND2X2 U1585 ( .A(A[11]), .B(n977), .Y(\ab[11][4] ) );
  AND2X2 U1586 ( .A(A[11]), .B(n978), .Y(\ab[11][3] ) );
  AND2X2 U1587 ( .A(A[11]), .B(n976), .Y(\ab[11][2] ) );
  AND2X2 U1588 ( .A(A[11]), .B(n980), .Y(\ab[11][1] ) );
  AND2X2 U1589 ( .A(A[11]), .B(n974), .Y(\ab[11][0] ) );
  AND2X2 U1590 ( .A(A[12]), .B(n1015), .Y(\ab[12][14] ) );
  NOR2X1 U1591 ( .A(A[11]), .B(n1051), .Y(\ab[11][15] ) );
  AND2X2 U1592 ( .A(A[12]), .B(n1013), .Y(\ab[12][13] ) );
  AND2X2 U1593 ( .A(A[12]), .B(n1011), .Y(\ab[12][12] ) );
  AND2X2 U1594 ( .A(A[12]), .B(n163), .Y(\ab[12][11] ) );
  AND2X2 U1595 ( .A(A[12]), .B(n1007), .Y(\ab[12][10] ) );
  AND2X2 U1596 ( .A(A[12]), .B(n507), .Y(\ab[12][9] ) );
  AND2X2 U1597 ( .A(A[12]), .B(n1005), .Y(\ab[12][8] ) );
  AND2X2 U1598 ( .A(A[12]), .B(n905), .Y(\ab[12][7] ) );
  AND2X2 U1599 ( .A(A[12]), .B(n969), .Y(\ab[12][6] ) );
  AND2X2 U1600 ( .A(A[12]), .B(n973), .Y(\ab[12][5] ) );
  AND2X2 U1601 ( .A(A[12]), .B(n977), .Y(\ab[12][4] ) );
  AND2X2 U1602 ( .A(A[12]), .B(n978), .Y(\ab[12][3] ) );
  AND2X2 U1603 ( .A(A[12]), .B(n976), .Y(\ab[12][2] ) );
  AND2X2 U1604 ( .A(A[12]), .B(n980), .Y(\ab[12][1] ) );
  AND2X2 U1605 ( .A(A[12]), .B(n974), .Y(\ab[12][0] ) );
  NOR2X1 U1606 ( .A(n1054), .B(n1037), .Y(\ab[13][14] ) );
  NOR2X1 U1607 ( .A(A[12]), .B(n1051), .Y(\ab[12][15] ) );
  NOR2X1 U1608 ( .A(n1054), .B(n1038), .Y(\ab[13][13] ) );
  NOR2X1 U1609 ( .A(n1054), .B(n1039), .Y(\ab[13][12] ) );
  NOR2X1 U1610 ( .A(n1054), .B(n1040), .Y(\ab[13][11] ) );
  NOR2X1 U1611 ( .A(n1054), .B(n1041), .Y(\ab[13][10] ) );
  NOR2X1 U1612 ( .A(n1054), .B(n1042), .Y(\ab[13][9] ) );
  NOR2X1 U1613 ( .A(n1054), .B(n1004), .Y(\ab[13][8] ) );
  NOR2X1 U1614 ( .A(n1054), .B(n1043), .Y(\ab[13][7] ) );
  NOR2X1 U1615 ( .A(n1054), .B(n1044), .Y(\ab[13][6] ) );
  NOR2X1 U1616 ( .A(n1054), .B(n1045), .Y(\ab[13][5] ) );
  NOR2X1 U1617 ( .A(n1054), .B(n1046), .Y(\ab[13][4] ) );
  NOR2X1 U1618 ( .A(n1054), .B(n1047), .Y(\ab[13][3] ) );
  NOR2X1 U1619 ( .A(n1054), .B(n1048), .Y(\ab[13][2] ) );
  NOR2X1 U1620 ( .A(n1054), .B(n1049), .Y(\ab[13][1] ) );
  NOR2X1 U1621 ( .A(n1054), .B(n989), .Y(\ab[13][0] ) );
  NOR2X1 U1622 ( .A(n1053), .B(n1037), .Y(\ab[14][14] ) );
  NOR2X1 U1623 ( .A(A[13]), .B(n1051), .Y(\ab[13][15] ) );
  NOR2X1 U1624 ( .A(n1053), .B(n1038), .Y(\ab[14][13] ) );
  NOR2X1 U1625 ( .A(n1053), .B(n1039), .Y(\ab[14][12] ) );
  NOR2X1 U1626 ( .A(n1053), .B(n1040), .Y(\ab[14][11] ) );
  NOR2X1 U1627 ( .A(n1053), .B(n1041), .Y(\ab[14][10] ) );
  NOR2X1 U1628 ( .A(n1053), .B(n1042), .Y(\ab[14][9] ) );
  NOR2X1 U1629 ( .A(n1053), .B(n1004), .Y(\ab[14][8] ) );
  NOR2X1 U1630 ( .A(n1053), .B(n1043), .Y(\ab[14][7] ) );
  NOR2X1 U1631 ( .A(n1053), .B(n1044), .Y(\ab[14][6] ) );
  NOR2X1 U1632 ( .A(n1053), .B(n1045), .Y(\ab[14][5] ) );
  NOR2X1 U1633 ( .A(n1053), .B(n1046), .Y(\ab[14][4] ) );
  NOR2X1 U1634 ( .A(n1053), .B(n1047), .Y(\ab[14][3] ) );
  NOR2X1 U1635 ( .A(n1053), .B(n1048), .Y(\ab[14][2] ) );
  NOR2X1 U1636 ( .A(n1053), .B(n1049), .Y(\ab[14][1] ) );
  NOR2X1 U1637 ( .A(n1053), .B(n989), .Y(\ab[14][0] ) );
  NOR2X1 U1638 ( .A(n1052), .B(n1051), .Y(\ab[15][15] ) );
  NOR2X1 U1639 ( .A(A[14]), .B(n1051), .Y(\ab[14][15] ) );
  AND2X2 U1640 ( .A(n974), .B(n402), .Y(PRODUCT[0]) );
  INVX2 U1641 ( .A(\CARRYB[15][15] ), .Y(n1050) );
  NOR2X1 U1642 ( .A(n507), .B(n1052), .Y(\ab[15][9] ) );
  NOR2X1 U1643 ( .A(n1005), .B(n1052), .Y(\ab[15][8] ) );
  NOR2X1 U1644 ( .A(n905), .B(n1052), .Y(\ab[15][7] ) );
  NOR2X1 U1645 ( .A(n969), .B(n1052), .Y(\ab[15][6] ) );
  NOR2X1 U1646 ( .A(n972), .B(n1052), .Y(\ab[15][5] ) );
  NOR2X1 U1647 ( .A(n977), .B(n1052), .Y(\ab[15][4] ) );
  NOR2X1 U1648 ( .A(n978), .B(n1052), .Y(\ab[15][3] ) );
  NOR2X1 U1649 ( .A(n976), .B(n1052), .Y(\ab[15][2] ) );
  NOR2X1 U1650 ( .A(n980), .B(n1052), .Y(\ab[15][1] ) );
  NOR2X1 U1651 ( .A(n1015), .B(n1052), .Y(\ab[15][14] ) );
  NOR2X1 U1652 ( .A(n1013), .B(n1052), .Y(\ab[15][13] ) );
  NOR2X1 U1653 ( .A(n1011), .B(n1052), .Y(\ab[15][12] ) );
  NOR2X1 U1654 ( .A(n163), .B(n1052), .Y(\ab[15][11] ) );
  NOR2X1 U1655 ( .A(n1007), .B(n1052), .Y(\ab[15][10] ) );
  NOR2X1 U1656 ( .A(n974), .B(n1052), .Y(\ab[15][0] ) );
endmodule


module matrix_math_DW01_add_23 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] ,
         \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64;
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2X2 U2 ( .A(n20), .B(n29), .Y(n2) );
  OR2X1 U3 ( .A(B[16]), .B(A[16]), .Y(n1) );
  OR2X1 U4 ( .A(A[16]), .B(B[16]), .Y(n54) );
  AND2X1 U5 ( .A(n29), .B(n30), .Y(n28) );
  INVX2 U6 ( .A(n44), .Y(n34) );
  INVX1 U7 ( .A(n31), .Y(n26) );
  NAND2X1 U8 ( .A(n3), .B(n2), .Y(n4) );
  NAND2X1 U9 ( .A(n4), .B(n35), .Y(n32) );
  INVX1 U10 ( .A(n34), .Y(n3) );
  INVX1 U11 ( .A(n27), .Y(n5) );
  INVX1 U12 ( .A(n5), .Y(n6) );
  INVX1 U13 ( .A(A[14]), .Y(n7) );
  INVX1 U14 ( .A(n7), .Y(n8) );
  OR2X1 U15 ( .A(n16), .B(n13), .Y(n60) );
  XNOR2X1 U16 ( .A(n50), .B(n9), .Y(SUM[18]) );
  NAND2X1 U17 ( .A(n40), .B(n45), .Y(n9) );
  INVX1 U18 ( .A(A[19]), .Y(n10) );
  INVX1 U19 ( .A(n10), .Y(n11) );
  OR2X2 U20 ( .A(A[15]), .B(B[15]), .Y(n12) );
  OR2X1 U21 ( .A(A[15]), .B(B[15]), .Y(n59) );
  INVX1 U22 ( .A(n41), .Y(n36) );
  BUFX2 U23 ( .A(B[14]), .Y(n13) );
  BUFX2 U24 ( .A(n1), .Y(n14) );
  AND2X2 U25 ( .A(n53), .B(n1), .Y(n15) );
  INVX1 U26 ( .A(n15), .Y(n46) );
  BUFX2 U27 ( .A(A[14]), .Y(n16) );
  XNOR2X1 U28 ( .A(n62), .B(n17), .Y(SUM[16]) );
  NAND2X1 U29 ( .A(n56), .B(n54), .Y(n17) );
  XOR2X1 U30 ( .A(n64), .B(n18), .Y(SUM[15]) );
  NAND2X1 U31 ( .A(n58), .B(n12), .Y(n18) );
  XNOR2X1 U32 ( .A(n55), .B(n19), .Y(SUM[17]) );
  AND2X2 U33 ( .A(n49), .B(n53), .Y(n19) );
  AND2X2 U34 ( .A(n15), .B(n45), .Y(n20) );
  XNOR2X1 U35 ( .A(n27), .B(n42), .Y(SUM[19]) );
  AND2X2 U36 ( .A(n64), .B(n60), .Y(SUM[14]) );
  NAND2X1 U37 ( .A(n57), .B(n58), .Y(n44) );
  NAND2X1 U38 ( .A(n58), .B(n63), .Y(n62) );
  XOR2X1 U39 ( .A(n22), .B(n23), .Y(SUM[21]) );
  XOR2X1 U40 ( .A(B[21]), .B(A[21]), .Y(n23) );
  NAND2X1 U41 ( .A(n24), .B(n25), .Y(n22) );
  OAI21X1 U42 ( .A(n26), .B(n6), .C(n28), .Y(n25) );
  XNOR2X1 U43 ( .A(n32), .B(n33), .Y(SUM[20]) );
  NAND2X1 U44 ( .A(n30), .B(n24), .Y(n33) );
  NAND2X1 U45 ( .A(B[20]), .B(A[20]), .Y(n24) );
  OR2X2 U46 ( .A(A[20]), .B(B[20]), .Y(n30) );
  AOI21X1 U47 ( .A(n36), .B(n29), .C(n37), .Y(n35) );
  NAND2X1 U48 ( .A(n31), .B(n38), .Y(n37) );
  NAND2X1 U49 ( .A(n39), .B(n29), .Y(n38) );
  INVX2 U50 ( .A(n40), .Y(n39) );
  NAND2X1 U51 ( .A(n31), .B(n29), .Y(n42) );
  OR2X2 U52 ( .A(A[19]), .B(B[19]), .Y(n29) );
  NAND2X1 U53 ( .A(n11), .B(B[19]), .Y(n31) );
  NAND3X1 U54 ( .A(n41), .B(n40), .C(n43), .Y(n27) );
  NAND2X1 U55 ( .A(n44), .B(n20), .Y(n43) );
  NAND2X1 U56 ( .A(n47), .B(n45), .Y(n41) );
  NAND2X1 U57 ( .A(n48), .B(n49), .Y(n47) );
  OR2X2 U58 ( .A(A[18]), .B(B[18]), .Y(n45) );
  NAND2X1 U59 ( .A(B[18]), .B(A[18]), .Y(n40) );
  OAI21X1 U60 ( .A(n34), .B(n46), .C(n51), .Y(n50) );
  AND2X2 U61 ( .A(n48), .B(n49), .Y(n51) );
  NAND2X1 U62 ( .A(n53), .B(n52), .Y(n48) );
  OR2X2 U63 ( .A(A[17]), .B(B[17]), .Y(n53) );
  NAND2X1 U64 ( .A(B[17]), .B(A[17]), .Y(n49) );
  AOI21X1 U65 ( .A(n44), .B(n14), .C(n52), .Y(n55) );
  INVX2 U66 ( .A(n56), .Y(n52) );
  NAND2X1 U67 ( .A(n12), .B(n61), .Y(n57) );
  AND2X2 U68 ( .A(A[14]), .B(B[14]), .Y(n61) );
  NAND2X1 U69 ( .A(A[16]), .B(B[16]), .Y(n56) );
  NAND2X1 U70 ( .A(n59), .B(n61), .Y(n63) );
  NAND2X1 U71 ( .A(A[15]), .B(B[15]), .Y(n58) );
  NAND2X1 U72 ( .A(n8), .B(n13), .Y(n64) );
endmodule


module matrix_math_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][15] ,
         \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][1] , \ab[1][0] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] ,
         \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][14] ,
         \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] ,
         \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] ,
         \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][13] , \SUMB[15][15] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[15][0] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , ZA, ZB,
         \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[21] , \A2[14] , n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign ZA = A[15];
  assign ZB = B[15];

  FAX1 S4_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .C(\SUMB[14][8] ), .YC(
        \CARRYB[15][7] ), .YS(\SUMB[15][7] ) );
  FAX1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .C(\SUMB[14][9] ), .YC(
        \CARRYB[15][8] ), .YS(\SUMB[15][8] ) );
  FAX1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .C(\SUMB[14][10] ), .YC(
        \CARRYB[15][9] ), .YS(\SUMB[15][9] ) );
  FAX1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .C(\SUMB[14][11] ), 
        .YC(\CARRYB[15][10] ), .YS(\SUMB[15][10] ) );
  FAX1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .C(\SUMB[14][12] ), 
        .YC(\CARRYB[15][11] ), .YS(\SUMB[15][11] ) );
  FAX1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .C(\SUMB[14][13] ), 
        .YC(\CARRYB[15][12] ), .YS(\SUMB[15][12] ) );
  FAX1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .C(\SUMB[14][14] ), 
        .YC(\CARRYB[15][13] ), .YS(\SUMB[15][13] ) );
  FAX1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .C(\ab[14][15] ), .YC(
        \CARRYB[15][14] ), .YS(\SUMB[15][14] ) );
  FAX1 S14_15 ( .A(n1096), .B(n1095), .C(\ab[15][15] ), .YC(\CARRYB[15][15] ), 
        .YS(\SUMB[15][15] ) );
  FAX1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .C(\SUMB[13][10] ), 
        .YC(\CARRYB[14][9] ), .YS(\SUMB[14][9] ) );
  FAX1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .C(\SUMB[13][11] ), 
        .YC(\CARRYB[14][10] ), .YS(\SUMB[14][10] ) );
  FAX1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .C(\SUMB[13][12] ), 
        .YC(\CARRYB[14][11] ), .YS(\SUMB[14][11] ) );
  FAX1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .C(\SUMB[13][13] ), 
        .YC(\CARRYB[14][12] ), .YS(\SUMB[14][12] ) );
  FAX1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .C(\SUMB[13][14] ), 
        .YC(\CARRYB[14][13] ), .YS(\SUMB[14][13] ) );
  FAX1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .C(\ab[13][15] ), 
        .YC(\CARRYB[14][14] ), .YS(\SUMB[14][14] ) );
  FAX1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .C(\SUMB[12][11] ), 
        .YC(\CARRYB[13][10] ), .YS(\SUMB[13][10] ) );
  FAX1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .C(\SUMB[12][12] ), 
        .YC(\CARRYB[13][11] ), .YS(\SUMB[13][11] ) );
  FAX1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .C(\SUMB[12][13] ), 
        .YC(\CARRYB[13][12] ), .YS(\SUMB[13][12] ) );
  FAX1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .C(\SUMB[12][14] ), 
        .YC(\CARRYB[13][13] ), .YS(\SUMB[13][13] ) );
  FAX1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .C(\ab[12][15] ), 
        .YC(\CARRYB[13][14] ), .YS(\SUMB[13][14] ) );
  FAX1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .C(\SUMB[11][9] ), .YC(
        \CARRYB[12][8] ), .YS(\SUMB[12][8] ) );
  FAX1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .C(\SUMB[11][11] ), 
        .YC(\CARRYB[12][10] ), .YS(\SUMB[12][10] ) );
  FAX1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .C(\SUMB[11][12] ), 
        .YC(\CARRYB[12][11] ), .YS(\SUMB[12][11] ) );
  FAX1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .C(\SUMB[11][13] ), 
        .YC(\CARRYB[12][12] ), .YS(\SUMB[12][12] ) );
  FAX1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .C(\SUMB[11][14] ), 
        .YC(\CARRYB[12][13] ), .YS(\SUMB[12][13] ) );
  FAX1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .C(\ab[11][15] ), 
        .YC(\CARRYB[12][14] ), .YS(\SUMB[12][14] ) );
  FAX1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .C(\SUMB[10][12] ), 
        .YC(\CARRYB[11][11] ), .YS(\SUMB[11][11] ) );
  FAX1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .C(\SUMB[10][13] ), 
        .YC(\CARRYB[11][12] ), .YS(\SUMB[11][12] ) );
  FAX1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .C(\SUMB[10][14] ), 
        .YC(\CARRYB[11][13] ), .YS(\SUMB[11][13] ) );
  FAX1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .C(\ab[10][15] ), 
        .YC(\CARRYB[11][14] ), .YS(\SUMB[11][14] ) );
  FAX1 S1_10_0 ( .A(\ab[10][0] ), .B(\SUMB[9][1] ), .C(\CARRYB[9][0] ), .YC(
        \CARRYB[10][0] ), .YS(\A1[8] ) );
  FAX1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .C(\SUMB[9][14] ), 
        .YC(\CARRYB[10][13] ), .YS(\SUMB[10][13] ) );
  FAX1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .C(\ab[9][15] ), .YC(
        \CARRYB[10][14] ), .YS(\SUMB[10][14] ) );
  FAX1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .C(\SUMB[8][2] ), .YC(
        \CARRYB[9][1] ), .YS(\SUMB[9][1] ) );
  FAX1 S2_9_11 ( .A(\CARRYB[8][11] ), .B(\ab[9][11] ), .C(\SUMB[8][12] ), .YC(
        \CARRYB[9][11] ), .YS(\SUMB[9][11] ) );
  FAX1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .C(\ab[8][15] ), .YC(
        \CARRYB[9][14] ), .YS(\SUMB[9][14] ) );
  FAX1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .C(\SUMB[7][13] ), .YC(
        \CARRYB[8][12] ), .YS(\SUMB[8][12] ) );
  FAX1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .C(\SUMB[7][14] ), .YC(
        \CARRYB[8][13] ), .YS(\SUMB[8][13] ) );
  FAX1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .C(\ab[7][15] ), .YC(
        \CARRYB[8][14] ), .YS(\SUMB[8][14] ) );
  FAX1 S2_7_11 ( .A(\ab[7][11] ), .B(n251), .C(\SUMB[6][12] ), .YC(
        \CARRYB[7][11] ), .YS(\SUMB[7][11] ) );
  FAX1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .C(\ab[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S1_6_0 ( .A(\CARRYB[5][0] ), .B(\ab[6][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S1_5_0 ( .A(\CARRYB[4][0] ), .B(\ab[5][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(\A1[3] ) );
  FAX1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .C(\ab[4][15] ), .YC(
        \CARRYB[5][14] ), .YS(\SUMB[5][14] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S3_3_14 ( .A(\ab[3][14] ), .B(\ab[2][15] ), .C(\CARRYB[2][14] ), .YC(
        \CARRYB[3][14] ), .YS(\SUMB[3][14] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n1020), .C(\SUMB[1][1] ), .YC(
        \CARRYB[2][0] ), .YS(\A1[0] ) );
  matrix_math_DW01_add_23 FS_1 ( .A({n1094, \A1[28] , \A1[27] , \A1[26] , 
        \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , 
        \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n95, n94, n93, n92, 
        n91, n90, n89, n88, \A2[21] , n1019, n1018, n1017, n1016, n1015, n1014, 
        \A2[14] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, PRODUCT[23:2]}) );
  AND2X2 U2 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(n3) );
  BUFX2 U3 ( .A(n739), .Y(n4) );
  NAND3X1 U4 ( .A(n670), .B(n669), .C(n668), .Y(n5) );
  BUFX2 U5 ( .A(n741), .Y(n6) );
  NAND3X1 U6 ( .A(n820), .B(n821), .C(n822), .Y(n7) );
  BUFX2 U7 ( .A(n603), .Y(n8) );
  XOR2X1 U8 ( .A(n62), .B(n9), .Y(\SUMB[3][11] ) );
  XNOR2X1 U9 ( .A(\CARRYB[2][11] ), .B(\ab[3][11] ), .Y(n9) );
  XNOR2X1 U10 ( .A(n10), .B(n11), .Y(\SUMB[6][4] ) );
  XOR2X1 U11 ( .A(\SUMB[5][5] ), .B(\ab[6][4] ), .Y(n10) );
  INVX1 U12 ( .A(\CARRYB[5][4] ), .Y(n11) );
  BUFX2 U13 ( .A(n187), .Y(n12) );
  XOR2X1 U14 ( .A(n13), .B(n36), .Y(\SUMB[13][1] ) );
  XOR2X1 U15 ( .A(\CARRYB[12][1] ), .B(n271), .Y(n13) );
  INVX1 U16 ( .A(\SUMB[12][2] ), .Y(n36) );
  INVX2 U17 ( .A(n913), .Y(n914) );
  XOR2X1 U18 ( .A(n14), .B(\ab[2][9] ), .Y(n15) );
  NAND2X1 U19 ( .A(\ab[0][10] ), .B(n429), .Y(n14) );
  XNOR2X1 U20 ( .A(n15), .B(\SUMB[1][10] ), .Y(\SUMB[2][9] ) );
  BUFX2 U21 ( .A(n896), .Y(n16) );
  BUFX2 U22 ( .A(\SUMB[5][2] ), .Y(n17) );
  XOR2X1 U23 ( .A(\CARRYB[9][5] ), .B(\ab[10][5] ), .Y(n281) );
  NAND2X1 U24 ( .A(\ab[8][3] ), .B(n141), .Y(n18) );
  XOR2X1 U25 ( .A(\CARRYB[11][4] ), .B(\ab[12][4] ), .Y(n47) );
  BUFX2 U26 ( .A(\SUMB[10][11] ), .Y(n19) );
  BUFX2 U27 ( .A(n188), .Y(n20) );
  XNOR2X1 U28 ( .A(n21), .B(n218), .Y(\SUMB[5][8] ) );
  XOR2X1 U29 ( .A(\CARRYB[4][8] ), .B(\ab[5][8] ), .Y(n21) );
  XNOR2X1 U30 ( .A(n22), .B(n45), .Y(\SUMB[7][7] ) );
  XOR2X1 U31 ( .A(\CARRYB[6][7] ), .B(\ab[7][7] ), .Y(n22) );
  XNOR2X1 U32 ( .A(\CARRYB[2][9] ), .B(n23), .Y(n182) );
  INVX8 U33 ( .A(\ab[3][9] ), .Y(n23) );
  BUFX2 U34 ( .A(n958), .Y(n24) );
  INVX2 U35 ( .A(\SUMB[4][5] ), .Y(n527) );
  INVX2 U36 ( .A(\SUMB[6][3] ), .Y(n453) );
  XNOR2X1 U37 ( .A(n25), .B(\SUMB[9][7] ), .Y(\SUMB[10][6] ) );
  XNOR2X1 U38 ( .A(\CARRYB[9][6] ), .B(\ab[10][6] ), .Y(n25) );
  XNOR2X1 U39 ( .A(n26), .B(\SUMB[6][9] ), .Y(\SUMB[7][8] ) );
  XNOR2X1 U40 ( .A(\CARRYB[6][8] ), .B(n40), .Y(n26) );
  BUFX2 U41 ( .A(n787), .Y(n27) );
  XNOR2X1 U42 ( .A(n235), .B(n179), .Y(n28) );
  XNOR2X1 U43 ( .A(n29), .B(\SUMB[9][5] ), .Y(\SUMB[10][4] ) );
  XNOR2X1 U44 ( .A(\CARRYB[9][4] ), .B(\ab[10][4] ), .Y(n29) );
  XNOR2X1 U45 ( .A(n30), .B(\SUMB[13][6] ), .Y(\SUMB[14][5] ) );
  XNOR2X1 U46 ( .A(\CARRYB[13][5] ), .B(n48), .Y(n30) );
  XOR2X1 U47 ( .A(n454), .B(n31), .Y(n227) );
  INVX8 U48 ( .A(\ab[12][3] ), .Y(n31) );
  BUFX2 U49 ( .A(\SUMB[12][1] ), .Y(n32) );
  XOR2X1 U50 ( .A(n394), .B(n33), .Y(n432) );
  INVX8 U51 ( .A(\ab[14][2] ), .Y(n33) );
  XOR2X1 U52 ( .A(\CARRYB[8][3] ), .B(n34), .Y(n724) );
  INVX8 U53 ( .A(\ab[9][3] ), .Y(n34) );
  XOR2X1 U54 ( .A(n35), .B(n76), .Y(\SUMB[9][5] ) );
  XOR2X1 U55 ( .A(\CARRYB[8][5] ), .B(\ab[9][5] ), .Y(n35) );
  XOR2X1 U56 ( .A(\CARRYB[11][5] ), .B(n37), .Y(n132) );
  INVX8 U57 ( .A(\ab[12][5] ), .Y(n37) );
  XOR2X1 U58 ( .A(n38), .B(\SUMB[4][8] ), .Y(\SUMB[5][7] ) );
  XOR2X1 U59 ( .A(\CARRYB[4][7] ), .B(\ab[5][7] ), .Y(n38) );
  BUFX2 U60 ( .A(n959), .Y(n39) );
  INVX8 U61 ( .A(n526), .Y(n40) );
  XNOR2X1 U62 ( .A(n41), .B(\SUMB[5][9] ), .Y(\SUMB[6][8] ) );
  XNOR2X1 U63 ( .A(\CARRYB[5][8] ), .B(\ab[6][8] ), .Y(n41) );
  BUFX2 U64 ( .A(A[1]), .Y(n42) );
  INVX1 U65 ( .A(A[1]), .Y(n430) );
  BUFX2 U66 ( .A(\SUMB[2][14] ), .Y(n43) );
  BUFX2 U67 ( .A(\SUMB[4][13] ), .Y(n44) );
  INVX2 U68 ( .A(\SUMB[4][9] ), .Y(n218) );
  INVX2 U69 ( .A(\SUMB[6][8] ), .Y(n45) );
  XOR2X1 U70 ( .A(n46), .B(\CARRYB[11][6] ), .Y(\SUMB[12][6] ) );
  XNOR2X1 U71 ( .A(\SUMB[11][7] ), .B(n355), .Y(n46) );
  XOR2X1 U72 ( .A(n47), .B(\SUMB[11][5] ), .Y(\SUMB[12][4] ) );
  INVX8 U73 ( .A(n397), .Y(n48) );
  XOR2X1 U74 ( .A(n49), .B(n511), .Y(\SUMB[2][14] ) );
  XNOR2X1 U75 ( .A(n196), .B(\ab[2][14] ), .Y(n49) );
  INVX4 U76 ( .A(B[13]), .Y(n1057) );
  XNOR2X1 U77 ( .A(n50), .B(\SUMB[1][13] ), .Y(\SUMB[2][12] ) );
  XNOR2X1 U78 ( .A(n388), .B(\ab[2][12] ), .Y(n50) );
  XNOR2X1 U79 ( .A(\CARRYB[14][3] ), .B(n80), .Y(n146) );
  BUFX2 U80 ( .A(n872), .Y(n51) );
  XNOR2X1 U81 ( .A(n835), .B(n52), .Y(n541) );
  INVX8 U82 ( .A(\ab[6][9] ), .Y(n52) );
  XNOR2X1 U83 ( .A(n53), .B(\SUMB[10][8] ), .Y(\SUMB[11][7] ) );
  XOR2X1 U84 ( .A(\CARRYB[10][7] ), .B(n654), .Y(n53) );
  XNOR2X1 U85 ( .A(n54), .B(\SUMB[14][6] ), .Y(\SUMB[15][5] ) );
  XNOR2X1 U86 ( .A(\CARRYB[14][5] ), .B(\ab[15][5] ), .Y(n54) );
  XOR2X1 U87 ( .A(n182), .B(n68), .Y(n55) );
  NAND3X1 U88 ( .A(n598), .B(n599), .C(n600), .Y(n56) );
  INVX2 U89 ( .A(\SUMB[12][4] ), .Y(n387) );
  BUFX2 U90 ( .A(n899), .Y(n57) );
  XNOR2X1 U91 ( .A(\CARRYB[7][6] ), .B(n58), .Y(n107) );
  INVX8 U92 ( .A(n224), .Y(n58) );
  INVX2 U93 ( .A(\SUMB[2][11] ), .Y(n59) );
  INVX2 U94 ( .A(n59), .Y(n60) );
  XOR2X1 U95 ( .A(n61), .B(\SUMB[1][12] ), .Y(\SUMB[2][11] ) );
  XNOR2X1 U96 ( .A(n174), .B(\ab[2][11] ), .Y(n61) );
  INVX1 U97 ( .A(\SUMB[2][12] ), .Y(n62) );
  XNOR2X1 U98 ( .A(\CARRYB[13][3] ), .B(n474), .Y(n63) );
  XOR2X1 U99 ( .A(n797), .B(n64), .Y(n386) );
  INVX8 U100 ( .A(n73), .Y(n64) );
  XOR2X1 U101 ( .A(n65), .B(\SUMB[4][10] ), .Y(\SUMB[5][9] ) );
  XNOR2X1 U102 ( .A(\CARRYB[4][9] ), .B(n173), .Y(n65) );
  INVX4 U103 ( .A(ZB), .Y(n1095) );
  XNOR2X1 U104 ( .A(n66), .B(\SUMB[5][13] ), .Y(\SUMB[6][12] ) );
  XNOR2X1 U105 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .Y(n66) );
  AND2X1 U106 ( .A(\SUMB[15][6] ), .B(\CARRYB[15][5] ), .Y(n1019) );
  XOR2X1 U107 ( .A(n67), .B(n276), .Y(\SUMB[12][1] ) );
  XOR2X1 U108 ( .A(n666), .B(\ab[12][1] ), .Y(n67) );
  XOR2X1 U109 ( .A(n216), .B(n272), .Y(n68) );
  AND2X2 U110 ( .A(\ab[0][10] ), .B(n429), .Y(n69) );
  XOR2X1 U111 ( .A(\CARRYB[10][4] ), .B(n70), .Y(n240) );
  INVX8 U112 ( .A(\ab[11][4] ), .Y(n70) );
  XOR2X1 U113 ( .A(\CARRYB[14][2] ), .B(n71), .Y(n255) );
  INVX8 U114 ( .A(n72), .Y(n71) );
  INVX8 U115 ( .A(\ab[15][2] ), .Y(n72) );
  INVX8 U116 ( .A(\ab[13][3] ), .Y(n73) );
  BUFX2 U117 ( .A(\SUMB[9][4] ), .Y(n74) );
  XOR2X1 U118 ( .A(\CARRYB[12][2] ), .B(n75), .Y(n164) );
  INVX8 U119 ( .A(\ab[13][2] ), .Y(n75) );
  XOR2X1 U120 ( .A(n107), .B(n217), .Y(n76) );
  XOR2X1 U121 ( .A(n123), .B(n121), .Y(n77) );
  INVX4 U122 ( .A(n1053), .Y(n1054) );
  INVX1 U123 ( .A(B[11]), .Y(n1053) );
  AND2X2 U124 ( .A(\ab[0][3] ), .B(n1022), .Y(n78) );
  AND2X2 U125 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n1021) );
  XOR2X1 U126 ( .A(\SUMB[7][9] ), .B(n79), .Y(n81) );
  INVX8 U127 ( .A(n211), .Y(n79) );
  INVX8 U128 ( .A(\ab[15][3] ), .Y(n80) );
  XOR2X1 U129 ( .A(n81), .B(\CARRYB[7][8] ), .Y(\SUMB[8][8] ) );
  XOR2X1 U130 ( .A(n181), .B(n356), .Y(n82) );
  XOR2X1 U131 ( .A(\SUMB[5][12] ), .B(\ab[6][11] ), .Y(n83) );
  XOR2X1 U132 ( .A(n83), .B(\CARRYB[5][11] ), .Y(\SUMB[6][11] ) );
  NAND2X1 U133 ( .A(\CARRYB[5][11] ), .B(\SUMB[5][12] ), .Y(n84) );
  NAND2X1 U134 ( .A(\CARRYB[5][11] ), .B(\ab[6][11] ), .Y(n85) );
  NAND2X1 U135 ( .A(\SUMB[5][12] ), .B(\ab[6][11] ), .Y(n86) );
  NAND3X1 U136 ( .A(n85), .B(n84), .C(n86), .Y(\CARRYB[6][11] ) );
  INVX2 U137 ( .A(\SUMB[7][6] ), .Y(n235) );
  XOR2X1 U138 ( .A(\CARRYB[5][7] ), .B(n87), .Y(n715) );
  INVX8 U139 ( .A(\ab[6][7] ), .Y(n87) );
  INVX2 U140 ( .A(\ab[10][7] ), .Y(n119) );
  INVX2 U141 ( .A(\ab[10][3] ), .Y(n577) );
  INVX2 U142 ( .A(\ab[5][9] ), .Y(n173) );
  INVX2 U143 ( .A(\ab[5][10] ), .Y(n213) );
  INVX2 U144 ( .A(\ab[5][6] ), .Y(n532) );
  INVX2 U145 ( .A(\ab[4][6] ), .Y(n208) );
  INVX2 U146 ( .A(\ab[8][8] ), .Y(n211) );
  INVX2 U147 ( .A(\ab[13][3] ), .Y(n520) );
  INVX2 U148 ( .A(\ab[12][6] ), .Y(n355) );
  INVX2 U149 ( .A(\ab[10][2] ), .Y(n731) );
  INVX2 U150 ( .A(\ab[12][2] ), .Y(n448) );
  INVX2 U151 ( .A(\ab[7][8] ), .Y(n526) );
  INVX2 U152 ( .A(\ab[7][9] ), .Y(n234) );
  INVX2 U153 ( .A(\ab[6][6] ), .Y(n228) );
  INVX2 U154 ( .A(\ab[6][5] ), .Y(n150) );
  INVX2 U155 ( .A(\ab[5][5] ), .Y(n434) );
  INVX2 U156 ( .A(\ab[8][6] ), .Y(n224) );
  INVX2 U157 ( .A(\ab[14][3] ), .Y(n474) );
  INVX2 U158 ( .A(\ab[13][4] ), .Y(n590) );
  INVX2 U159 ( .A(\ab[8][2] ), .Y(n463) );
  INVX2 U160 ( .A(n1034), .Y(n1035) );
  INVX2 U161 ( .A(\ab[14][5] ), .Y(n397) );
  INVX2 U162 ( .A(\ab[15][6] ), .Y(n540) );
  INVX2 U163 ( .A(n1080), .Y(n1081) );
  INVX2 U164 ( .A(\ab[13][1] ), .Y(n271) );
  INVX2 U165 ( .A(\ab[11][10] ), .Y(n197) );
  INVX2 U166 ( .A(n1046), .Y(n1047) );
  AND2X2 U167 ( .A(\SUMB[15][8] ), .B(\CARRYB[15][7] ), .Y(n88) );
  AND2X2 U168 ( .A(\SUMB[15][9] ), .B(\CARRYB[15][8] ), .Y(n89) );
  AND2X2 U169 ( .A(\SUMB[15][10] ), .B(\CARRYB[15][9] ), .Y(n90) );
  AND2X2 U170 ( .A(\SUMB[15][11] ), .B(\CARRYB[15][10] ), .Y(n91) );
  AND2X2 U171 ( .A(\SUMB[15][12] ), .B(\CARRYB[15][11] ), .Y(n92) );
  AND2X2 U172 ( .A(\SUMB[15][13] ), .B(\CARRYB[15][12] ), .Y(n93) );
  AND2X2 U173 ( .A(\SUMB[15][14] ), .B(\CARRYB[15][13] ), .Y(n94) );
  AND2X2 U174 ( .A(\SUMB[15][15] ), .B(\CARRYB[15][14] ), .Y(n95) );
  AND2X2 U175 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n96) );
  AND2X2 U176 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n97) );
  INVX2 U177 ( .A(n169), .Y(n104) );
  AND2X1 U178 ( .A(n789), .B(n791), .Y(n98) );
  AND2X1 U179 ( .A(n381), .B(n380), .Y(n99) );
  INVX2 U180 ( .A(\ab[11][3] ), .Y(n464) );
  BUFX2 U181 ( .A(\SUMB[4][7] ), .Y(n100) );
  BUFX2 U182 ( .A(\SUMB[5][6] ), .Y(n101) );
  XOR2X1 U183 ( .A(\SUMB[3][11] ), .B(n102), .Y(\SUMB[4][10] ) );
  XOR2X1 U184 ( .A(\CARRYB[3][10] ), .B(\ab[4][10] ), .Y(n102) );
  INVX2 U185 ( .A(n1061), .Y(n103) );
  INVX4 U186 ( .A(n1061), .Y(n1062) );
  INVX1 U187 ( .A(\SUMB[11][2] ), .Y(n276) );
  INVX2 U188 ( .A(\ab[2][10] ), .Y(n169) );
  INVX1 U189 ( .A(n1061), .Y(n105) );
  BUFX2 U190 ( .A(\ab[2][11] ), .Y(n106) );
  XOR2X1 U191 ( .A(n107), .B(n217), .Y(\SUMB[8][6] ) );
  INVX1 U192 ( .A(\SUMB[10][3] ), .Y(n149) );
  AND2X2 U193 ( .A(n42), .B(n1045), .Y(\ab[1][6] ) );
  AND2X1 U194 ( .A(n983), .B(B[1]), .Y(\ab[1][1] ) );
  NAND3X1 U195 ( .A(n368), .B(n367), .C(n369), .Y(n108) );
  NAND3X1 U196 ( .A(n881), .B(n882), .C(n883), .Y(n109) );
  BUFX2 U197 ( .A(n845), .Y(n110) );
  NAND3X1 U198 ( .A(n496), .B(n497), .C(n498), .Y(n111) );
  XNOR2X1 U199 ( .A(n112), .B(\SUMB[10][4] ), .Y(\SUMB[11][3] ) );
  XNOR2X1 U200 ( .A(n1028), .B(n464), .Y(n112) );
  AND2X1 U201 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(n186) );
  BUFX2 U202 ( .A(\SUMB[15][0] ), .Y(n113) );
  INVX1 U203 ( .A(\CARRYB[15][0] ), .Y(n114) );
  INVX1 U204 ( .A(n114), .Y(n115) );
  NAND3X1 U205 ( .A(n12), .B(n20), .C(n189), .Y(n116) );
  BUFX2 U206 ( .A(n873), .Y(n117) );
  XOR2X1 U207 ( .A(n118), .B(\SUMB[5][7] ), .Y(\SUMB[6][6] ) );
  XNOR2X1 U208 ( .A(\CARRYB[5][6] ), .B(n228), .Y(n118) );
  XOR2X1 U209 ( .A(\CARRYB[9][7] ), .B(n119), .Y(n273) );
  XOR2X1 U210 ( .A(n255), .B(n183), .Y(\SUMB[15][2] ) );
  NAND3X1 U211 ( .A(n385), .B(n384), .C(n383), .Y(\CARRYB[2][11] ) );
  XNOR2X1 U212 ( .A(n1025), .B(\ab[2][13] ), .Y(n779) );
  NAND3X1 U213 ( .A(n554), .B(n556), .C(n555), .Y(n394) );
  BUFX2 U214 ( .A(n846), .Y(n120) );
  XNOR2X1 U215 ( .A(n164), .B(n200), .Y(n121) );
  XOR2X1 U216 ( .A(n589), .B(n122), .Y(\SUMB[8][4] ) );
  XNOR2X1 U217 ( .A(\CARRYB[7][4] ), .B(\ab[8][4] ), .Y(n122) );
  XOR2X1 U218 ( .A(n123), .B(n121), .Y(\SUMB[14][1] ) );
  XNOR2X1 U219 ( .A(n1030), .B(\ab[14][1] ), .Y(n123) );
  NAND3X1 U220 ( .A(n716), .B(n717), .C(n718), .Y(n124) );
  NAND3X1 U221 ( .A(n844), .B(n110), .C(n120), .Y(n125) );
  XOR2X1 U222 ( .A(n724), .B(n329), .Y(n126) );
  XNOR2X1 U223 ( .A(n127), .B(n28), .Y(\SUMB[9][4] ) );
  XNOR2X1 U224 ( .A(\CARRYB[8][4] ), .B(\ab[9][4] ), .Y(n127) );
  NAND3X1 U225 ( .A(n823), .B(n824), .C(n825), .Y(n128) );
  NAND3X1 U226 ( .A(n891), .B(n892), .C(n893), .Y(n129) );
  NAND3X1 U227 ( .A(n338), .B(n337), .C(n339), .Y(n130) );
  BUFX2 U228 ( .A(n751), .Y(n131) );
  XNOR2X1 U229 ( .A(n132), .B(\SUMB[11][6] ), .Y(\SUMB[12][5] ) );
  XNOR2X1 U230 ( .A(n133), .B(\SUMB[10][7] ), .Y(\SUMB[11][6] ) );
  XNOR2X1 U231 ( .A(\CARRYB[10][6] ), .B(\ab[11][6] ), .Y(n133) );
  NAND3X1 U232 ( .A(n535), .B(n533), .C(n534), .Y(n134) );
  NAND3X1 U233 ( .A(n331), .B(n332), .C(n333), .Y(n135) );
  NAND3X1 U234 ( .A(n743), .B(n744), .C(n745), .Y(n136) );
  XOR2X1 U235 ( .A(n432), .B(n433), .Y(n137) );
  NAND3X1 U236 ( .A(n515), .B(n516), .C(n517), .Y(n138) );
  BUFX2 U237 ( .A(\CARRYB[15][2] ), .Y(n139) );
  NAND3X1 U238 ( .A(n606), .B(n605), .C(n607), .Y(n140) );
  NAND3X1 U239 ( .A(n725), .B(n727), .C(n726), .Y(n141) );
  NAND3X1 U240 ( .A(n598), .B(n599), .C(n600), .Y(n142) );
  NAND3X1 U241 ( .A(n904), .B(n906), .C(n905), .Y(n143) );
  NAND3X1 U242 ( .A(n635), .B(n637), .C(n636), .Y(n144) );
  NAND3X1 U243 ( .A(n989), .B(n990), .C(n991), .Y(n145) );
  XOR2X1 U244 ( .A(n146), .B(\SUMB[14][4] ), .Y(\SUMB[15][3] ) );
  XOR2X1 U245 ( .A(n147), .B(n575), .Y(\SUMB[7][4] ) );
  XOR2X1 U246 ( .A(\CARRYB[6][4] ), .B(\ab[7][4] ), .Y(n147) );
  XOR2X1 U247 ( .A(n545), .B(\ab[11][2] ), .Y(n148) );
  XNOR2X1 U248 ( .A(n148), .B(n149), .Y(\SUMB[11][2] ) );
  XOR2X1 U249 ( .A(\CARRYB[5][5] ), .B(n150), .Y(n167) );
  XOR2X1 U250 ( .A(\CARRYB[14][1] ), .B(\ab[15][1] ), .Y(n547) );
  XNOR2X1 U251 ( .A(n151), .B(\SUMB[8][8] ), .Y(\SUMB[9][7] ) );
  XNOR2X1 U252 ( .A(\CARRYB[8][7] ), .B(\ab[9][7] ), .Y(n151) );
  XOR2X1 U253 ( .A(n152), .B(\SUMB[6][6] ), .Y(\SUMB[7][5] ) );
  XOR2X1 U254 ( .A(\CARRYB[6][5] ), .B(\ab[7][5] ), .Y(n152) );
  BUFX2 U255 ( .A(n1065), .Y(n153) );
  XOR2X1 U256 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .Y(n154) );
  XOR2X1 U257 ( .A(n154), .B(\SUMB[12][10] ), .Y(\SUMB[13][9] ) );
  XOR2X1 U258 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .Y(n155) );
  XOR2X1 U259 ( .A(n155), .B(\SUMB[13][9] ), .Y(\SUMB[14][8] ) );
  NAND2X1 U260 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .Y(n156) );
  NAND2X1 U261 ( .A(\ab[13][9] ), .B(\SUMB[12][10] ), .Y(n157) );
  NAND2X1 U262 ( .A(\CARRYB[12][9] ), .B(\SUMB[12][10] ), .Y(n158) );
  NAND3X1 U263 ( .A(n156), .B(n157), .C(n158), .Y(\CARRYB[13][9] ) );
  NAND2X1 U264 ( .A(\ab[14][8] ), .B(n108), .Y(n159) );
  NAND2X1 U265 ( .A(\ab[14][8] ), .B(\SUMB[13][9] ), .Y(n160) );
  NAND2X1 U266 ( .A(n108), .B(\SUMB[13][9] ), .Y(n161) );
  NAND3X1 U267 ( .A(n159), .B(n160), .C(n161), .Y(\CARRYB[14][8] ) );
  BUFX2 U268 ( .A(\SUMB[3][13] ), .Y(n162) );
  NAND3X1 U269 ( .A(n782), .B(n780), .C(n781), .Y(n163) );
  XNOR2X1 U270 ( .A(n164), .B(n200), .Y(\SUMB[13][2] ) );
  BUFX2 U271 ( .A(\CARRYB[4][7] ), .Y(n165) );
  XNOR2X1 U272 ( .A(n166), .B(\ab[1][8] ), .Y(\SUMB[1][8] ) );
  NAND2X1 U273 ( .A(B[9]), .B(n1062), .Y(n166) );
  XNOR2X1 U274 ( .A(n167), .B(n101), .Y(\SUMB[6][5] ) );
  INVX1 U275 ( .A(\SUMB[3][7] ), .Y(n254) );
  XNOR2X1 U276 ( .A(n168), .B(n314), .Y(\SUMB[4][9] ) );
  XOR2X1 U277 ( .A(\CARRYB[3][9] ), .B(\ab[4][9] ), .Y(n168) );
  BUFX2 U278 ( .A(n466), .Y(n170) );
  XNOR2X1 U279 ( .A(\CARRYB[9][8] ), .B(\ab[10][8] ), .Y(n357) );
  INVX2 U280 ( .A(\SUMB[2][13] ), .Y(n356) );
  INVX2 U281 ( .A(\CARRYB[3][7] ), .Y(n947) );
  XNOR2X1 U282 ( .A(n171), .B(n74), .Y(\SUMB[10][3] ) );
  XOR2X1 U283 ( .A(\CARRYB[9][3] ), .B(n577), .Y(n171) );
  XNOR2X1 U284 ( .A(n172), .B(\SUMB[8][10] ), .Y(\SUMB[9][9] ) );
  XNOR2X1 U285 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .Y(n172) );
  INVX2 U286 ( .A(n430), .Y(n252) );
  NAND2X1 U287 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(n174) );
  XOR2X1 U288 ( .A(ZA), .B(ZB), .Y(n175) );
  XOR2X1 U289 ( .A(n113), .B(n175), .Y(\A1[13] ) );
  NAND2X1 U290 ( .A(\SUMB[15][0] ), .B(ZA), .Y(n176) );
  NAND2X1 U291 ( .A(\SUMB[15][0] ), .B(ZB), .Y(n177) );
  NAND2X1 U292 ( .A(ZA), .B(ZB), .Y(n178) );
  NAND3X1 U293 ( .A(n178), .B(n177), .C(n176), .Y(\A2[14] ) );
  NAND2X1 U294 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .Y(n928) );
  AND2X1 U295 ( .A(\SUMB[15][4] ), .B(\CARRYB[15][3] ), .Y(n1017) );
  XNOR2X1 U296 ( .A(n235), .B(n179), .Y(\SUMB[8][5] ) );
  XOR2X1 U297 ( .A(\CARRYB[7][5] ), .B(\ab[8][5] ), .Y(n179) );
  XOR2X1 U298 ( .A(\SUMB[12][8] ), .B(n180), .Y(\SUMB[13][7] ) );
  XOR2X1 U299 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .Y(n180) );
  XOR2X1 U300 ( .A(n181), .B(n356), .Y(\SUMB[3][12] ) );
  XNOR2X1 U301 ( .A(\CARRYB[2][12] ), .B(\ab[3][12] ), .Y(n181) );
  INVX2 U302 ( .A(\SUMB[13][3] ), .Y(n433) );
  XOR2X1 U303 ( .A(n182), .B(n68), .Y(\SUMB[3][9] ) );
  NAND2X1 U304 ( .A(n260), .B(n261), .Y(n183) );
  NAND3X1 U305 ( .A(n384), .B(n383), .C(n385), .Y(n184) );
  AND2X2 U306 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(n185) );
  NAND2X1 U307 ( .A(\SUMB[1][13] ), .B(n388), .Y(n187) );
  NAND2X1 U308 ( .A(\SUMB[1][13] ), .B(\ab[2][12] ), .Y(n188) );
  NAND2X1 U309 ( .A(n388), .B(\ab[2][12] ), .Y(n189) );
  NAND3X1 U310 ( .A(n189), .B(n187), .C(n188), .Y(\CARRYB[2][12] ) );
  XNOR2X1 U311 ( .A(n190), .B(\SUMB[4][12] ), .Y(\SUMB[5][11] ) );
  XOR2X1 U312 ( .A(n831), .B(\ab[5][11] ), .Y(n190) );
  XOR2X1 U313 ( .A(\ab[4][14] ), .B(\ab[3][15] ), .Y(n191) );
  XOR2X1 U314 ( .A(\CARRYB[3][14] ), .B(n191), .Y(\SUMB[4][14] ) );
  NAND2X1 U315 ( .A(\CARRYB[3][14] ), .B(\ab[4][14] ), .Y(n192) );
  NAND2X1 U316 ( .A(\CARRYB[3][14] ), .B(\ab[3][15] ), .Y(n193) );
  NAND2X1 U317 ( .A(\ab[4][14] ), .B(\ab[3][15] ), .Y(n194) );
  NAND3X1 U318 ( .A(n193), .B(n192), .C(n194), .Y(\CARRYB[4][14] ) );
  AND2X2 U319 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Y(n195) );
  AND2X2 U320 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Y(n196) );
  XNOR2X1 U321 ( .A(n197), .B(\SUMB[10][11] ), .Y(n374) );
  XOR2X1 U322 ( .A(\SUMB[15][7] ), .B(\CARRYB[15][6] ), .Y(\A1[20] ) );
  NAND2X1 U323 ( .A(\ab[4][10] ), .B(n834), .Y(n198) );
  INVX2 U324 ( .A(n833), .Y(n834) );
  XNOR2X1 U325 ( .A(n199), .B(\SUMB[9][12] ), .Y(\SUMB[10][11] ) );
  XNOR2X1 U326 ( .A(\CARRYB[9][11] ), .B(\ab[10][11] ), .Y(n199) );
  XOR2X1 U327 ( .A(n227), .B(n431), .Y(n200) );
  NAND3X1 U328 ( .A(n786), .B(n788), .C(n27), .Y(n201) );
  INVX2 U329 ( .A(\SUMB[11][4] ), .Y(n431) );
  XNOR2X1 U330 ( .A(n202), .B(\SUMB[3][8] ), .Y(\SUMB[4][7] ) );
  XNOR2X1 U331 ( .A(n947), .B(n680), .Y(n202) );
  NAND2X1 U332 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .Y(n203) );
  BUFX2 U333 ( .A(n865), .Y(n204) );
  BUFX2 U334 ( .A(\SUMB[2][2] ), .Y(n205) );
  NAND2X1 U335 ( .A(n447), .B(n446), .Y(n206) );
  XNOR2X1 U336 ( .A(n207), .B(\SUMB[2][9] ), .Y(\SUMB[3][8] ) );
  XNOR2X1 U337 ( .A(\CARRYB[2][8] ), .B(\ab[3][8] ), .Y(n207) );
  INVX2 U338 ( .A(\SUMB[7][7] ), .Y(n217) );
  XNOR2X1 U339 ( .A(n208), .B(n138), .Y(n212) );
  XOR2X1 U340 ( .A(n225), .B(n209), .Y(\SUMB[10][9] ) );
  INVX2 U341 ( .A(\SUMB[9][10] ), .Y(n209) );
  AND2X2 U342 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n210) );
  XNOR2X1 U343 ( .A(n212), .B(n254), .Y(\SUMB[4][6] ) );
  XOR2X1 U344 ( .A(\CARRYB[14][4] ), .B(\ab[15][4] ), .Y(n309) );
  XOR2X1 U345 ( .A(\CARRYB[4][10] ), .B(n213), .Y(n214) );
  XNOR2X1 U346 ( .A(n214), .B(n267), .Y(\SUMB[5][10] ) );
  XOR2X1 U347 ( .A(n215), .B(n222), .Y(\SUMB[3][6] ) );
  XNOR2X1 U348 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .Y(n215) );
  XOR2X1 U349 ( .A(n216), .B(n272), .Y(\SUMB[2][10] ) );
  INVX1 U350 ( .A(\SUMB[1][11] ), .Y(n216) );
  NAND3X1 U351 ( .A(n499), .B(n500), .C(n501), .Y(n219) );
  NAND3X1 U352 ( .A(n817), .B(n818), .C(n819), .Y(n220) );
  NAND3X1 U353 ( .A(n644), .B(n646), .C(n645), .Y(n221) );
  INVX1 U354 ( .A(\SUMB[2][7] ), .Y(n222) );
  XNOR2X1 U355 ( .A(n976), .B(n223), .Y(\SUMB[2][6] ) );
  INVX1 U356 ( .A(\SUMB[1][7] ), .Y(n223) );
  XNOR2X1 U357 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .Y(n225) );
  XNOR2X1 U358 ( .A(n226), .B(\SUMB[8][11] ), .Y(\SUMB[9][10] ) );
  XNOR2X1 U359 ( .A(\CARRYB[8][10] ), .B(\ab[9][10] ), .Y(n226) );
  XOR2X1 U360 ( .A(n227), .B(n431), .Y(\SUMB[12][3] ) );
  NAND3X1 U361 ( .A(n884), .B(n885), .C(n886), .Y(n229) );
  AND2X1 U362 ( .A(\SUMB[15][5] ), .B(\CARRYB[15][4] ), .Y(n1018) );
  XNOR2X1 U363 ( .A(n274), .B(n230), .Y(\SUMB[3][7] ) );
  XOR2X1 U364 ( .A(\CARRYB[2][7] ), .B(\ab[3][7] ), .Y(n230) );
  BUFX4 U365 ( .A(\SUMB[6][5] ), .Y(n575) );
  BUFX2 U366 ( .A(\CARRYB[10][5] ), .Y(n231) );
  NAND3X1 U367 ( .A(n461), .B(n462), .C(n460), .Y(n232) );
  XOR2X1 U368 ( .A(n233), .B(n55), .Y(\SUMB[4][8] ) );
  XNOR2X1 U369 ( .A(n913), .B(\ab[4][8] ), .Y(n233) );
  XOR2X1 U370 ( .A(\CARRYB[6][9] ), .B(n234), .Y(n421) );
  NAND2X1 U371 ( .A(\ab[10][1] ), .B(n1026), .Y(n236) );
  BUFX2 U372 ( .A(\SUMB[3][5] ), .Y(n237) );
  XNOR2X1 U373 ( .A(\ab[5][12] ), .B(n829), .Y(n503) );
  INVX2 U374 ( .A(n829), .Y(n830) );
  NAND3X1 U375 ( .A(n868), .B(n870), .C(n869), .Y(n238) );
  XNOR2X1 U376 ( .A(n239), .B(\SUMB[2][6] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U377 ( .A(\ab[3][5] ), .B(n985), .Y(n239) );
  XOR2X1 U378 ( .A(n240), .B(n241), .Y(\SUMB[11][4] ) );
  XOR2X1 U379 ( .A(n281), .B(n519), .Y(n241) );
  NAND2X1 U380 ( .A(n790), .B(n98), .Y(n946) );
  BUFX2 U381 ( .A(n750), .Y(n242) );
  INVX1 U382 ( .A(\CARRYB[4][2] ), .Y(n573) );
  INVX1 U383 ( .A(\ab[3][13] ), .Y(n244) );
  XNOR2X1 U384 ( .A(n243), .B(\SUMB[7][11] ), .Y(\SUMB[8][10] ) );
  XNOR2X1 U385 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .Y(n243) );
  XNOR2X1 U386 ( .A(n244), .B(\CARRYB[2][13] ), .Y(n874) );
  INVX2 U387 ( .A(\SUMB[8][4] ), .Y(n329) );
  BUFX2 U388 ( .A(\SUMB[15][3] ), .Y(n245) );
  XNOR2X1 U389 ( .A(n246), .B(\SUMB[14][7] ), .Y(\SUMB[15][6] ) );
  XOR2X1 U390 ( .A(\CARRYB[14][6] ), .B(n540), .Y(n246) );
  NAND2X1 U391 ( .A(n379), .B(n99), .Y(n594) );
  INVX2 U392 ( .A(\CARRYB[11][1] ), .Y(n666) );
  XNOR2X1 U393 ( .A(n247), .B(\SUMB[10][10] ), .Y(\SUMB[11][9] ) );
  XNOR2X1 U394 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .Y(n247) );
  XOR2X1 U395 ( .A(n248), .B(n527), .Y(\SUMB[5][4] ) );
  XNOR2X1 U396 ( .A(\CARRYB[4][4] ), .B(\ab[5][4] ), .Y(n248) );
  INVX1 U397 ( .A(B[7]), .Y(n1046) );
  XNOR2X1 U398 ( .A(n249), .B(n722), .Y(\SUMB[2][8] ) );
  XOR2X1 U399 ( .A(\ab[2][8] ), .B(n440), .Y(n249) );
  INVX2 U400 ( .A(\CARRYB[6][11] ), .Y(n250) );
  INVX4 U401 ( .A(n250), .Y(n251) );
  XNOR2X1 U402 ( .A(n253), .B(n262), .Y(\SUMB[2][7] ) );
  XOR2X1 U403 ( .A(\ab[2][7] ), .B(n270), .Y(n253) );
  INVX1 U404 ( .A(n839), .Y(n840) );
  INVX2 U405 ( .A(\CARRYB[15][0] ), .Y(n749) );
  NAND2X1 U406 ( .A(\SUMB[14][3] ), .B(n201), .Y(n256) );
  NAND2X1 U407 ( .A(\SUMB[14][3] ), .B(\ab[15][2] ), .Y(n257) );
  NAND2X1 U408 ( .A(n201), .B(\ab[15][2] ), .Y(n258) );
  NAND3X1 U409 ( .A(n258), .B(n256), .C(n257), .Y(\CARRYB[15][2] ) );
  NAND2X1 U410 ( .A(\SUMB[13][4] ), .B(n277), .Y(n260) );
  NAND2X1 U411 ( .A(n63), .B(n259), .Y(n261) );
  NAND2X1 U412 ( .A(n260), .B(n261), .Y(\SUMB[14][3] ) );
  INVX1 U413 ( .A(\SUMB[13][4] ), .Y(n259) );
  BUFX2 U414 ( .A(\SUMB[1][8] ), .Y(n262) );
  NAND3X1 U415 ( .A(n895), .B(n897), .C(n16), .Y(n263) );
  BUFX2 U416 ( .A(\SUMB[9][2] ), .Y(n264) );
  NAND3X1 U417 ( .A(n795), .B(n796), .C(n794), .Y(n265) );
  NAND3X1 U418 ( .A(n951), .B(n952), .C(n953), .Y(n266) );
  BUFX2 U419 ( .A(\SUMB[4][11] ), .Y(n267) );
  NAND3X1 U420 ( .A(n811), .B(n812), .C(n813), .Y(n268) );
  NAND3X1 U421 ( .A(n647), .B(n648), .C(n649), .Y(n269) );
  NAND2X1 U422 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(n270) );
  INVX1 U423 ( .A(n985), .Y(n986) );
  XOR2X1 U424 ( .A(n1024), .B(\ab[2][10] ), .Y(n272) );
  INVX1 U425 ( .A(\CARRYB[6][9] ), .Y(n839) );
  XNOR2X1 U426 ( .A(n273), .B(\SUMB[9][8] ), .Y(\SUMB[10][7] ) );
  INVX1 U427 ( .A(\SUMB[2][8] ), .Y(n274) );
  XNOR2X1 U428 ( .A(n956), .B(n275), .Y(\SUMB[9][6] ) );
  INVX1 U429 ( .A(\SUMB[8][7] ), .Y(n275) );
  XOR2X1 U430 ( .A(n678), .B(n474), .Y(n277) );
  BUFX2 U431 ( .A(\SUMB[3][6] ), .Y(n278) );
  BUFX2 U432 ( .A(\SUMB[10][2] ), .Y(n279) );
  INVX2 U433 ( .A(\SUMB[3][10] ), .Y(n314) );
  BUFX2 U434 ( .A(n740), .Y(n280) );
  XNOR2X1 U435 ( .A(n281), .B(n519), .Y(\SUMB[10][5] ) );
  XOR2X1 U436 ( .A(\CARRYB[6][13] ), .B(\ab[7][13] ), .Y(n282) );
  XOR2X1 U437 ( .A(n282), .B(\SUMB[6][14] ), .Y(\SUMB[7][13] ) );
  NAND2X1 U438 ( .A(\SUMB[6][14] ), .B(\CARRYB[6][13] ), .Y(n283) );
  NAND2X1 U439 ( .A(\SUMB[6][14] ), .B(\ab[7][13] ), .Y(n284) );
  NAND2X1 U440 ( .A(\CARRYB[6][13] ), .B(\ab[7][13] ), .Y(n285) );
  NAND3X1 U441 ( .A(n284), .B(n283), .C(n285), .Y(\CARRYB[7][13] ) );
  XOR2X1 U442 ( .A(\ab[5][15] ), .B(\ab[6][14] ), .Y(n286) );
  XOR2X1 U443 ( .A(\CARRYB[5][14] ), .B(n286), .Y(\SUMB[6][14] ) );
  NAND2X1 U444 ( .A(\CARRYB[5][14] ), .B(\ab[5][15] ), .Y(n287) );
  NAND2X1 U445 ( .A(\CARRYB[5][14] ), .B(\ab[6][14] ), .Y(n288) );
  NAND2X1 U446 ( .A(\ab[5][15] ), .B(\ab[6][14] ), .Y(n289) );
  NAND3X1 U447 ( .A(n288), .B(n287), .C(n289), .Y(\CARRYB[6][14] ) );
  XOR2X1 U448 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .Y(n290) );
  XOR2X1 U449 ( .A(n290), .B(\SUMB[8][14] ), .Y(\SUMB[9][13] ) );
  XOR2X1 U450 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .Y(n291) );
  XOR2X1 U451 ( .A(n291), .B(\SUMB[9][13] ), .Y(\SUMB[10][12] ) );
  NAND2X1 U452 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .Y(n292) );
  NAND2X1 U453 ( .A(\ab[9][13] ), .B(\SUMB[8][14] ), .Y(n293) );
  NAND2X1 U454 ( .A(\CARRYB[8][13] ), .B(\SUMB[8][14] ), .Y(n294) );
  NAND3X1 U455 ( .A(n292), .B(n293), .C(n294), .Y(\CARRYB[9][13] ) );
  NAND2X1 U456 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .Y(n295) );
  NAND2X1 U457 ( .A(\ab[10][12] ), .B(\SUMB[9][13] ), .Y(n296) );
  NAND2X1 U458 ( .A(\CARRYB[9][12] ), .B(\SUMB[9][13] ), .Y(n297) );
  NAND3X1 U459 ( .A(n295), .B(n296), .C(n297), .Y(\CARRYB[10][12] ) );
  BUFX2 U460 ( .A(A[0]), .Y(n298) );
  XOR2X1 U461 ( .A(\SUMB[1][5] ), .B(\ab[2][4] ), .Y(n299) );
  XOR2X1 U462 ( .A(n97), .B(n299), .Y(\SUMB[2][4] ) );
  NAND2X1 U463 ( .A(\SUMB[1][5] ), .B(n97), .Y(n300) );
  NAND2X1 U464 ( .A(n97), .B(\ab[2][4] ), .Y(n301) );
  NAND2X1 U465 ( .A(\SUMB[1][5] ), .B(\ab[2][4] ), .Y(n302) );
  NAND3X1 U466 ( .A(n301), .B(n300), .C(n302), .Y(\CARRYB[2][4] ) );
  BUFX2 U467 ( .A(\SUMB[4][3] ), .Y(n303) );
  INVX4 U468 ( .A(A[3]), .Y(n1066) );
  NAND2X1 U469 ( .A(\SUMB[4][10] ), .B(\CARRYB[4][9] ), .Y(n304) );
  NAND2X1 U470 ( .A(\SUMB[4][10] ), .B(\ab[5][9] ), .Y(n305) );
  NAND2X1 U471 ( .A(\CARRYB[4][9] ), .B(\ab[5][9] ), .Y(n306) );
  NAND3X1 U472 ( .A(n306), .B(n305), .C(n304), .Y(\CARRYB[5][9] ) );
  NAND3X1 U473 ( .A(n871), .B(n51), .C(n117), .Y(n307) );
  NAND3X1 U474 ( .A(n131), .B(n242), .C(n752), .Y(n308) );
  XOR2X1 U475 ( .A(n309), .B(\SUMB[14][5] ), .Y(\SUMB[15][4] ) );
  NAND2X1 U476 ( .A(\SUMB[14][5] ), .B(n129), .Y(n310) );
  NAND2X1 U477 ( .A(\SUMB[14][5] ), .B(\ab[15][4] ), .Y(n311) );
  NAND2X1 U478 ( .A(n129), .B(\ab[15][4] ), .Y(n312) );
  NAND3X1 U479 ( .A(n311), .B(n310), .C(n312), .Y(\CARRYB[15][4] ) );
  NAND3X1 U480 ( .A(n805), .B(n806), .C(n807), .Y(n313) );
  XNOR2X1 U481 ( .A(n315), .B(n126), .Y(\SUMB[10][2] ) );
  XOR2X1 U482 ( .A(\CARRYB[9][2] ), .B(n731), .Y(n315) );
  NAND3X1 U483 ( .A(n847), .B(n848), .C(n849), .Y(n316) );
  NAND3X1 U484 ( .A(n933), .B(n931), .C(n932), .Y(n317) );
  NAND3X1 U485 ( .A(n915), .B(n916), .C(n917), .Y(n318) );
  XOR2X1 U486 ( .A(n677), .B(n319), .Y(\SUMB[9][2] ) );
  INVX1 U487 ( .A(\SUMB[8][3] ), .Y(n319) );
  INVX1 U488 ( .A(\CARRYB[3][10] ), .Y(n833) );
  XNOR2X1 U489 ( .A(n320), .B(n136), .Y(\SUMB[13][4] ) );
  XOR2X1 U490 ( .A(\SUMB[12][5] ), .B(n590), .Y(n320) );
  AND2X2 U491 ( .A(n139), .B(n245), .Y(n1016) );
  NAND3X1 U492 ( .A(n965), .B(n963), .C(n964), .Y(n321) );
  NAND3X1 U493 ( .A(n856), .B(n858), .C(n857), .Y(n322) );
  NAND3X1 U494 ( .A(n583), .B(n584), .C(n582), .Y(n323) );
  NAND3X1 U495 ( .A(n706), .B(n708), .C(n707), .Y(n324) );
  NAND3X1 U496 ( .A(n198), .B(n816), .C(n815), .Y(n325) );
  NAND3X1 U497 ( .A(n888), .B(n890), .C(n889), .Y(n326) );
  NAND3X1 U498 ( .A(n808), .B(n809), .C(n810), .Y(n327) );
  NAND3X1 U499 ( .A(n465), .B(n170), .C(n467), .Y(n328) );
  XOR2X1 U500 ( .A(n724), .B(n329), .Y(\SUMB[9][3] ) );
  XOR2X1 U501 ( .A(\CARRYB[10][8] ), .B(\ab[11][8] ), .Y(n330) );
  XOR2X1 U502 ( .A(n330), .B(\SUMB[10][9] ), .Y(\SUMB[11][8] ) );
  NAND2X1 U503 ( .A(\ab[10][9] ), .B(n219), .Y(n331) );
  NAND2X1 U504 ( .A(\SUMB[9][10] ), .B(\ab[10][9] ), .Y(n332) );
  NAND2X1 U505 ( .A(n219), .B(\SUMB[9][10] ), .Y(n333) );
  NAND3X1 U506 ( .A(n331), .B(n332), .C(n333), .Y(\CARRYB[10][9] ) );
  NAND2X1 U507 ( .A(\ab[11][8] ), .B(n109), .Y(n334) );
  NAND2X1 U508 ( .A(\SUMB[10][9] ), .B(\ab[11][8] ), .Y(n335) );
  NAND2X1 U509 ( .A(n109), .B(\SUMB[10][9] ), .Y(n336) );
  NAND3X1 U510 ( .A(n334), .B(n335), .C(n336), .Y(\CARRYB[11][8] ) );
  INVX2 U511 ( .A(\CARRYB[15][5] ), .Y(n510) );
  NAND2X1 U512 ( .A(\SUMB[7][7] ), .B(n143), .Y(n337) );
  NAND2X1 U513 ( .A(\SUMB[7][7] ), .B(\ab[8][6] ), .Y(n338) );
  NAND2X1 U514 ( .A(n143), .B(\ab[8][6] ), .Y(n339) );
  NAND3X1 U515 ( .A(n338), .B(n337), .C(n339), .Y(\CARRYB[8][6] ) );
  NAND3X1 U516 ( .A(n4), .B(n280), .C(n6), .Y(n340) );
  NAND3X1 U517 ( .A(n559), .B(n558), .C(n557), .Y(n341) );
  INVX2 U518 ( .A(n831), .Y(n832) );
  XOR2X1 U519 ( .A(\SUMB[10][1] ), .B(\ab[11][0] ), .Y(n342) );
  XOR2X1 U520 ( .A(\CARRYB[10][0] ), .B(n342), .Y(\A1[9] ) );
  NAND2X1 U521 ( .A(\CARRYB[10][0] ), .B(\SUMB[10][1] ), .Y(n343) );
  NAND2X1 U522 ( .A(\CARRYB[10][0] ), .B(\ab[11][0] ), .Y(n344) );
  NAND2X1 U523 ( .A(\SUMB[10][1] ), .B(\ab[11][0] ), .Y(n345) );
  NAND3X1 U524 ( .A(n344), .B(n343), .C(n345), .Y(\CARRYB[11][0] ) );
  INVX1 U525 ( .A(\CARRYB[11][0] ), .Y(n866) );
  XNOR2X1 U526 ( .A(n346), .B(\SUMB[6][11] ), .Y(\SUMB[7][10] ) );
  XNOR2X1 U527 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .Y(n346) );
  INVX2 U528 ( .A(n866), .Y(n867) );
  NAND3X1 U529 ( .A(n236), .B(n720), .C(n721), .Y(n347) );
  INVX1 U530 ( .A(n524), .Y(n348) );
  NAND3X1 U531 ( .A(n977), .B(n978), .C(n979), .Y(n349) );
  INVX1 U532 ( .A(\SUMB[4][4] ), .Y(n522) );
  NAND2X1 U533 ( .A(\SUMB[4][11] ), .B(n325), .Y(n350) );
  NAND2X1 U534 ( .A(\SUMB[4][11] ), .B(\ab[5][10] ), .Y(n351) );
  NAND2X1 U535 ( .A(n325), .B(\ab[5][10] ), .Y(n352) );
  NAND3X1 U536 ( .A(n351), .B(n350), .C(n352), .Y(\CARRYB[5][10] ) );
  XOR2X1 U537 ( .A(n354), .B(n353), .Y(\SUMB[6][3] ) );
  XNOR2X1 U538 ( .A(n142), .B(\ab[6][3] ), .Y(n353) );
  INVX1 U539 ( .A(\SUMB[5][4] ), .Y(n354) );
  XNOR2X1 U540 ( .A(n426), .B(n264), .Y(\SUMB[10][1] ) );
  INVX1 U541 ( .A(n1056), .Y(n1084) );
  XNOR2X1 U542 ( .A(n357), .B(\SUMB[9][9] ), .Y(\SUMB[10][8] ) );
  XOR2X1 U543 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .Y(n358) );
  XOR2X1 U544 ( .A(n358), .B(\SUMB[5][14] ), .Y(\SUMB[6][13] ) );
  XOR2X1 U545 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .Y(n359) );
  XOR2X1 U546 ( .A(n359), .B(\SUMB[6][13] ), .Y(\SUMB[7][12] ) );
  NAND2X1 U547 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .Y(n360) );
  NAND2X1 U548 ( .A(\ab[6][13] ), .B(\SUMB[5][14] ), .Y(n361) );
  NAND2X1 U549 ( .A(\CARRYB[5][13] ), .B(\SUMB[5][14] ), .Y(n362) );
  NAND3X1 U550 ( .A(n360), .B(n361), .C(n362), .Y(\CARRYB[6][13] ) );
  NAND2X1 U551 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .Y(n363) );
  NAND2X1 U552 ( .A(\ab[7][12] ), .B(\SUMB[6][13] ), .Y(n364) );
  NAND2X1 U553 ( .A(\CARRYB[6][12] ), .B(\SUMB[6][13] ), .Y(n365) );
  NAND3X1 U554 ( .A(n363), .B(n364), .C(n365), .Y(\CARRYB[7][12] ) );
  XOR2X1 U555 ( .A(\CARRYB[12][8] ), .B(\ab[13][8] ), .Y(n366) );
  XOR2X1 U556 ( .A(\SUMB[12][9] ), .B(n366), .Y(\SUMB[13][8] ) );
  NAND2X1 U557 ( .A(\SUMB[12][9] ), .B(\CARRYB[12][8] ), .Y(n367) );
  NAND2X1 U558 ( .A(\SUMB[12][9] ), .B(\ab[13][8] ), .Y(n368) );
  NAND2X1 U559 ( .A(\CARRYB[12][8] ), .B(\ab[13][8] ), .Y(n369) );
  NAND3X1 U560 ( .A(n368), .B(n367), .C(n369), .Y(\CARRYB[13][8] ) );
  XOR2X1 U561 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .Y(n370) );
  XOR2X1 U562 ( .A(n370), .B(\SUMB[9][11] ), .Y(\SUMB[10][10] ) );
  NAND2X1 U563 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .Y(n371) );
  NAND2X1 U564 ( .A(\ab[10][10] ), .B(\SUMB[9][11] ), .Y(n372) );
  NAND2X1 U565 ( .A(\CARRYB[9][10] ), .B(\SUMB[9][11] ), .Y(n373) );
  NAND3X1 U566 ( .A(n371), .B(n372), .C(n373), .Y(\CARRYB[10][10] ) );
  XOR2X1 U567 ( .A(n374), .B(\CARRYB[10][10] ), .Y(\SUMB[11][10] ) );
  NAND2X1 U568 ( .A(\ab[11][10] ), .B(n19), .Y(n375) );
  NAND2X1 U569 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .Y(n376) );
  NAND2X1 U570 ( .A(n19), .B(\CARRYB[10][10] ), .Y(n377) );
  NAND3X1 U571 ( .A(n375), .B(n376), .C(n377), .Y(\CARRYB[11][10] ) );
  XNOR2X1 U572 ( .A(n435), .B(\SUMB[8][9] ), .Y(\SUMB[9][8] ) );
  XOR2X1 U573 ( .A(n347), .B(\ab[11][1] ), .Y(n378) );
  XOR2X1 U574 ( .A(n279), .B(n378), .Y(\SUMB[11][1] ) );
  NAND2X1 U575 ( .A(\CARRYB[10][1] ), .B(\SUMB[10][2] ), .Y(n379) );
  NAND2X1 U576 ( .A(\SUMB[10][2] ), .B(\ab[11][1] ), .Y(n380) );
  NAND2X1 U577 ( .A(\CARRYB[10][1] ), .B(\ab[11][1] ), .Y(n381) );
  NAND3X1 U578 ( .A(n380), .B(n379), .C(n381), .Y(\CARRYB[11][1] ) );
  INVX1 U579 ( .A(n1045), .Y(n1088) );
  XNOR2X1 U580 ( .A(n382), .B(\SUMB[4][6] ), .Y(\SUMB[5][5] ) );
  XOR2X1 U581 ( .A(\CARRYB[4][5] ), .B(n434), .Y(n382) );
  NAND2X1 U582 ( .A(\SUMB[1][12] ), .B(n186), .Y(n383) );
  NAND2X1 U583 ( .A(\SUMB[1][12] ), .B(n106), .Y(n384) );
  NAND2X1 U584 ( .A(n186), .B(n106), .Y(n385) );
  INVX4 U585 ( .A(B[12]), .Y(n1055) );
  XOR2X1 U586 ( .A(n386), .B(n387), .Y(\SUMB[13][3] ) );
  AND2X2 U587 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Y(n388) );
  NAND3X1 U588 ( .A(n709), .B(n710), .C(n711), .Y(n389) );
  NAND3X1 U589 ( .A(n457), .B(n456), .C(n458), .Y(n390) );
  NAND3X1 U590 ( .A(n512), .B(n513), .C(n514), .Y(n391) );
  XNOR2X1 U591 ( .A(\ab[0][10] ), .B(n392), .Y(\SUMB[1][9] ) );
  NAND2X1 U592 ( .A(n983), .B(n1050), .Y(n392) );
  NAND3X1 U593 ( .A(n565), .B(n563), .C(n564), .Y(n393) );
  NAND3X1 U594 ( .A(n898), .B(n900), .C(n57), .Y(n395) );
  NAND3X1 U595 ( .A(n934), .B(n935), .C(n936), .Y(n396) );
  INVX1 U596 ( .A(\CARRYB[10][7] ), .Y(n657) );
  XOR2X1 U597 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .Y(n398) );
  XOR2X1 U598 ( .A(n398), .B(\SUMB[8][13] ), .Y(\SUMB[9][12] ) );
  NAND2X1 U599 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .Y(n399) );
  NAND2X1 U600 ( .A(\ab[9][12] ), .B(\SUMB[8][13] ), .Y(n400) );
  NAND2X1 U601 ( .A(\CARRYB[8][12] ), .B(\SUMB[8][13] ), .Y(n401) );
  NAND3X1 U602 ( .A(n399), .B(n400), .C(n401), .Y(\CARRYB[9][12] ) );
  NAND2X1 U603 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .Y(n402) );
  NAND2X1 U604 ( .A(\ab[10][11] ), .B(\SUMB[9][12] ), .Y(n403) );
  NAND2X1 U605 ( .A(\CARRYB[9][11] ), .B(\SUMB[9][12] ), .Y(n404) );
  NAND3X1 U606 ( .A(n402), .B(n403), .C(n404), .Y(\CARRYB[10][11] ) );
  XOR2X1 U607 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .Y(n405) );
  XOR2X1 U608 ( .A(n405), .B(\SUMB[4][14] ), .Y(\SUMB[5][13] ) );
  NAND2X1 U609 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .Y(n406) );
  NAND2X1 U610 ( .A(\ab[5][13] ), .B(\SUMB[4][14] ), .Y(n407) );
  NAND2X1 U611 ( .A(\CARRYB[4][13] ), .B(\SUMB[4][14] ), .Y(n408) );
  NAND3X1 U612 ( .A(n406), .B(n407), .C(n408), .Y(\CARRYB[5][13] ) );
  NAND2X1 U613 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .Y(n409) );
  NAND2X1 U614 ( .A(\ab[6][12] ), .B(\SUMB[5][13] ), .Y(n410) );
  NAND2X1 U615 ( .A(\CARRYB[5][12] ), .B(\SUMB[5][13] ), .Y(n411) );
  NAND3X1 U616 ( .A(n409), .B(n410), .C(n411), .Y(\CARRYB[6][12] ) );
  XNOR2X1 U617 ( .A(n412), .B(\SUMB[5][11] ), .Y(\SUMB[6][10] ) );
  XOR2X1 U618 ( .A(\ab[6][10] ), .B(n837), .Y(n412) );
  XOR2X1 U619 ( .A(\SUMB[11][1] ), .B(\ab[12][0] ), .Y(n413) );
  XOR2X1 U620 ( .A(n867), .B(n413), .Y(\A1[10] ) );
  NAND2X1 U621 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Y(n414) );
  NAND2X1 U622 ( .A(\CARRYB[11][0] ), .B(\ab[12][0] ), .Y(n415) );
  NAND2X1 U623 ( .A(\SUMB[11][1] ), .B(\ab[12][0] ), .Y(n416) );
  NAND3X1 U624 ( .A(n415), .B(n416), .C(n414), .Y(\CARRYB[12][0] ) );
  BUFX2 U625 ( .A(\SUMB[5][3] ), .Y(n417) );
  NAND3X1 U626 ( .A(n864), .B(n863), .C(n204), .Y(n418) );
  NAND3X1 U627 ( .A(n980), .B(n982), .C(n981), .Y(n419) );
  NAND3X1 U628 ( .A(n472), .B(n471), .C(n473), .Y(n420) );
  XNOR2X1 U629 ( .A(n421), .B(\SUMB[6][10] ), .Y(\SUMB[7][9] ) );
  NAND3X1 U630 ( .A(n960), .B(n961), .C(n962), .Y(n422) );
  NAND2X1 U631 ( .A(\ab[7][2] ), .B(n5), .Y(n423) );
  BUFX2 U632 ( .A(\SUMB[2][5] ), .Y(n424) );
  XOR2X1 U633 ( .A(n425), .B(n660), .Y(\SUMB[2][5] ) );
  XNOR2X1 U634 ( .A(n439), .B(\ab[2][5] ), .Y(n425) );
  XNOR2X1 U635 ( .A(n1026), .B(\ab[10][1] ), .Y(n426) );
  NAND3X1 U636 ( .A(n203), .B(n638), .C(n639), .Y(n427) );
  NAND3X1 U637 ( .A(n998), .B(n997), .C(n999), .Y(n428) );
  AND2X2 U638 ( .A(n983), .B(n1050), .Y(n429) );
  INVX2 U639 ( .A(A[1]), .Y(n1063) );
  AND2X2 U640 ( .A(n252), .B(B[8]), .Y(\ab[1][8] ) );
  XOR2X1 U641 ( .A(n432), .B(n433), .Y(\SUMB[14][2] ) );
  INVX1 U642 ( .A(\SUMB[7][5] ), .Y(n589) );
  INVX2 U643 ( .A(\ab[1][15] ), .Y(n511) );
  XNOR2X1 U644 ( .A(\CARRYB[8][8] ), .B(\ab[9][8] ), .Y(n435) );
  NAND3X1 U645 ( .A(n630), .B(n631), .C(n632), .Y(n436) );
  AND2X2 U646 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(n437) );
  AND2X2 U647 ( .A(B[7]), .B(n983), .Y(\ab[1][7] ) );
  INVX1 U648 ( .A(\SUMB[1][6] ), .Y(n660) );
  INVX2 U649 ( .A(B[8]), .Y(n1048) );
  INVX2 U650 ( .A(n1063), .Y(n984) );
  BUFX2 U651 ( .A(\SUMB[3][4] ), .Y(n438) );
  AND2X2 U652 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n439) );
  AND2X2 U653 ( .A(n984), .B(B[2]), .Y(n1022) );
  AND2X2 U654 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(n440) );
  XNOR2X1 U655 ( .A(n420), .B(\ab[7][4] ), .Y(n441) );
  NAND3X1 U656 ( .A(n923), .B(n922), .C(n921), .Y(n442) );
  XNOR2X1 U657 ( .A(n443), .B(n424), .Y(\SUMB[3][4] ) );
  XOR2X1 U658 ( .A(n701), .B(\ab[3][4] ), .Y(n443) );
  NAND2X1 U659 ( .A(\SUMB[6][7] ), .B(n626), .Y(n446) );
  NAND2X1 U660 ( .A(n444), .B(n445), .Y(n447) );
  NAND2X1 U661 ( .A(n446), .B(n447), .Y(\SUMB[7][6] ) );
  INVX1 U662 ( .A(n626), .Y(n444) );
  INVX1 U663 ( .A(\SUMB[6][7] ), .Y(n445) );
  XNOR2X1 U664 ( .A(\CARRYB[11][2] ), .B(n448), .Y(n702) );
  XOR2X1 U665 ( .A(n449), .B(n450), .Y(\SUMB[1][7] ) );
  NAND2X1 U666 ( .A(n984), .B(B[7]), .Y(n449) );
  OR2X2 U667 ( .A(n1048), .B(n1061), .Y(n450) );
  INVX2 U668 ( .A(\CARRYB[7][3] ), .Y(n524) );
  INVX2 U669 ( .A(n1030), .Y(n1031) );
  AND2X2 U670 ( .A(ZB), .B(n1061), .Y(\ab[0][15] ) );
  NAND3X1 U671 ( .A(n712), .B(n713), .C(n714), .Y(n451) );
  XNOR2X1 U672 ( .A(n452), .B(\SUMB[13][8] ), .Y(\SUMB[14][7] ) );
  XNOR2X1 U673 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .Y(n452) );
  XNOR2X1 U674 ( .A(n1008), .B(n453), .Y(\SUMB[7][2] ) );
  NAND3X1 U675 ( .A(n703), .B(n704), .C(n705), .Y(n454) );
  NAND3X1 U676 ( .A(n907), .B(n908), .C(n909), .Y(n455) );
  NAND2X1 U677 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(n456) );
  NAND2X1 U678 ( .A(\CARRYB[7][8] ), .B(\ab[8][8] ), .Y(n457) );
  NAND2X1 U679 ( .A(\SUMB[7][9] ), .B(\ab[8][8] ), .Y(n458) );
  NAND3X1 U680 ( .A(n457), .B(n456), .C(n458), .Y(\CARRYB[8][8] ) );
  XOR2X1 U681 ( .A(\SUMB[10][6] ), .B(\ab[11][5] ), .Y(n459) );
  XOR2X1 U682 ( .A(n459), .B(n231), .Y(\SUMB[11][5] ) );
  NAND2X1 U683 ( .A(\SUMB[10][6] ), .B(\CARRYB[10][5] ), .Y(n460) );
  NAND2X1 U684 ( .A(\CARRYB[10][5] ), .B(\ab[11][5] ), .Y(n461) );
  NAND2X1 U685 ( .A(\SUMB[10][6] ), .B(\ab[11][5] ), .Y(n462) );
  NAND3X1 U686 ( .A(n461), .B(n462), .C(n460), .Y(\CARRYB[11][5] ) );
  XOR2X1 U687 ( .A(\CARRYB[7][2] ), .B(n463), .Y(n673) );
  INVX1 U688 ( .A(n1028), .Y(n1029) );
  NAND2X1 U689 ( .A(\ab[9][8] ), .B(n390), .Y(n465) );
  NAND2X1 U690 ( .A(\ab[9][8] ), .B(\SUMB[8][9] ), .Y(n466) );
  NAND2X1 U691 ( .A(\SUMB[8][9] ), .B(n390), .Y(n467) );
  NAND3X1 U692 ( .A(n465), .B(n466), .C(n467), .Y(\CARRYB[9][8] ) );
  NAND2X1 U693 ( .A(\ab[10][7] ), .B(n238), .Y(n468) );
  NAND2X1 U694 ( .A(\ab[10][7] ), .B(\SUMB[9][8] ), .Y(n469) );
  NAND2X1 U695 ( .A(n238), .B(\SUMB[9][8] ), .Y(n470) );
  NAND3X1 U696 ( .A(n468), .B(n469), .C(n470), .Y(\CARRYB[10][7] ) );
  AND2X2 U697 ( .A(B[9]), .B(n298), .Y(\ab[0][9] ) );
  NAND2X1 U698 ( .A(\SUMB[5][5] ), .B(\CARRYB[5][4] ), .Y(n471) );
  NAND2X1 U699 ( .A(\CARRYB[5][4] ), .B(\ab[6][4] ), .Y(n472) );
  NAND2X1 U700 ( .A(\SUMB[5][5] ), .B(\ab[6][4] ), .Y(n473) );
  NAND3X1 U701 ( .A(n472), .B(n473), .C(n471), .Y(\CARRYB[6][4] ) );
  XOR2X1 U702 ( .A(n475), .B(n278), .Y(\SUMB[4][5] ) );
  XOR2X1 U703 ( .A(\CARRYB[3][5] ), .B(\ab[4][5] ), .Y(n475) );
  BUFX2 U704 ( .A(\SUMB[3][3] ), .Y(n476) );
  XNOR2X1 U705 ( .A(n987), .B(n477), .Y(\SUMB[3][3] ) );
  INVX1 U706 ( .A(\SUMB[2][4] ), .Y(n477) );
  XNOR2X1 U707 ( .A(n676), .B(n478), .Y(\SUMB[7][3] ) );
  XOR2X1 U708 ( .A(\CARRYB[6][3] ), .B(\ab[7][3] ), .Y(n478) );
  XOR2X1 U709 ( .A(\SUMB[8][1] ), .B(\ab[9][0] ), .Y(n479) );
  XOR2X1 U710 ( .A(n479), .B(\CARRYB[8][0] ), .Y(\A1[7] ) );
  NAND2X1 U711 ( .A(\CARRYB[8][0] ), .B(\SUMB[8][1] ), .Y(n480) );
  NAND2X1 U712 ( .A(\CARRYB[8][0] ), .B(\ab[9][0] ), .Y(n481) );
  NAND2X1 U713 ( .A(\SUMB[8][1] ), .B(\ab[9][0] ), .Y(n482) );
  NAND3X1 U714 ( .A(n482), .B(n480), .C(n481), .Y(\CARRYB[9][0] ) );
  XOR2X1 U715 ( .A(\ab[2][1] ), .B(n96), .Y(n483) );
  XOR2X1 U716 ( .A(n483), .B(\SUMB[1][2] ), .Y(\SUMB[2][1] ) );
  XOR2X1 U717 ( .A(\CARRYB[2][0] ), .B(\ab[3][0] ), .Y(n484) );
  XOR2X1 U718 ( .A(n484), .B(\SUMB[2][1] ), .Y(\A1[1] ) );
  NAND2X1 U719 ( .A(\ab[2][1] ), .B(n96), .Y(n485) );
  NAND2X1 U720 ( .A(\ab[2][1] ), .B(\SUMB[1][2] ), .Y(n486) );
  NAND2X1 U721 ( .A(n96), .B(\SUMB[1][2] ), .Y(n487) );
  NAND3X1 U722 ( .A(n485), .B(n486), .C(n487), .Y(\CARRYB[2][1] ) );
  NAND2X1 U723 ( .A(\CARRYB[2][0] ), .B(\ab[3][0] ), .Y(n488) );
  NAND2X1 U724 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n489) );
  NAND2X1 U725 ( .A(\ab[3][0] ), .B(\SUMB[2][1] ), .Y(n490) );
  NAND3X1 U726 ( .A(n488), .B(n489), .C(n490), .Y(\CARRYB[3][0] ) );
  INVX1 U727 ( .A(n1037), .Y(n1092) );
  INVX2 U728 ( .A(\SUMB[9][6] ), .Y(n519) );
  NAND2X1 U729 ( .A(\SUMB[14][4] ), .B(n308), .Y(n491) );
  NAND2X1 U730 ( .A(\SUMB[14][4] ), .B(\ab[15][3] ), .Y(n492) );
  NAND2X1 U731 ( .A(n308), .B(\ab[15][3] ), .Y(n493) );
  NAND3X1 U732 ( .A(n492), .B(n491), .C(n493), .Y(\CARRYB[15][3] ) );
  NAND3X1 U733 ( .A(n957), .B(n39), .C(n24), .Y(n494) );
  NAND3X1 U734 ( .A(n746), .B(n748), .C(n747), .Y(n495) );
  NAND2X1 U735 ( .A(\ab[8][10] ), .B(n220), .Y(n496) );
  NAND2X1 U736 ( .A(\ab[8][10] ), .B(\SUMB[7][11] ), .Y(n497) );
  NAND2X1 U737 ( .A(n220), .B(\SUMB[7][11] ), .Y(n498) );
  NAND3X1 U738 ( .A(n496), .B(n497), .C(n498), .Y(\CARRYB[8][10] ) );
  NAND2X1 U739 ( .A(\ab[9][9] ), .B(n7), .Y(n499) );
  NAND2X1 U740 ( .A(\SUMB[8][10] ), .B(\ab[9][9] ), .Y(n500) );
  NAND2X1 U741 ( .A(n7), .B(\SUMB[8][10] ), .Y(n501) );
  NAND3X1 U742 ( .A(n499), .B(n500), .C(n501), .Y(\CARRYB[9][9] ) );
  XOR2X1 U743 ( .A(\CARRYB[3][13] ), .B(\ab[4][13] ), .Y(n502) );
  XOR2X1 U744 ( .A(n502), .B(\SUMB[3][14] ), .Y(\SUMB[4][13] ) );
  XOR2X1 U745 ( .A(n503), .B(n44), .Y(\SUMB[5][12] ) );
  NAND2X1 U746 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .Y(n504) );
  NAND2X1 U747 ( .A(\ab[4][13] ), .B(\SUMB[3][14] ), .Y(n505) );
  NAND2X1 U748 ( .A(\CARRYB[3][13] ), .B(\SUMB[3][14] ), .Y(n506) );
  NAND3X1 U749 ( .A(n504), .B(n505), .C(n506), .Y(\CARRYB[4][13] ) );
  NAND2X1 U750 ( .A(\ab[5][12] ), .B(n830), .Y(n507) );
  NAND2X1 U751 ( .A(\ab[5][12] ), .B(\SUMB[4][13] ), .Y(n508) );
  NAND2X1 U752 ( .A(n830), .B(\SUMB[4][13] ), .Y(n509) );
  NAND3X1 U753 ( .A(n507), .B(n508), .C(n509), .Y(\CARRYB[5][12] ) );
  XNOR2X1 U754 ( .A(\SUMB[15][6] ), .B(n510), .Y(\A1[19] ) );
  NAND2X1 U755 ( .A(\ab[2][7] ), .B(n437), .Y(n512) );
  NAND2X1 U756 ( .A(n437), .B(\SUMB[1][8] ), .Y(n513) );
  NAND2X1 U757 ( .A(\ab[2][7] ), .B(\SUMB[1][8] ), .Y(n514) );
  NAND3X1 U758 ( .A(n512), .B(n513), .C(n514), .Y(\CARRYB[2][7] ) );
  NAND2X1 U759 ( .A(\ab[3][6] ), .B(n349), .Y(n515) );
  NAND2X1 U760 ( .A(\ab[3][6] ), .B(\SUMB[2][7] ), .Y(n516) );
  NAND2X1 U761 ( .A(\SUMB[2][7] ), .B(n349), .Y(n517) );
  NAND3X1 U762 ( .A(n515), .B(n516), .C(n517), .Y(\CARRYB[3][6] ) );
  XNOR2X1 U763 ( .A(n441), .B(n575), .Y(n518) );
  XNOR2X1 U764 ( .A(n954), .B(n77), .Y(\SUMB[15][0] ) );
  OR2X2 U765 ( .A(n520), .B(n797), .Y(n783) );
  INVX1 U766 ( .A(n797), .Y(n798) );
  INVX1 U767 ( .A(n1060), .Y(n1082) );
  XOR2X1 U768 ( .A(n522), .B(n521), .Y(\SUMB[5][3] ) );
  XNOR2X1 U769 ( .A(n531), .B(\ab[5][3] ), .Y(n521) );
  NAND2X1 U770 ( .A(n523), .B(n524), .Y(n525) );
  NAND2X1 U771 ( .A(n973), .B(n525), .Y(n528) );
  INVX1 U772 ( .A(\ab[8][3] ), .Y(n523) );
  INVX2 U773 ( .A(n835), .Y(n836) );
  XNOR2X1 U774 ( .A(n528), .B(n518), .Y(\SUMB[8][3] ) );
  INVX4 U775 ( .A(n1048), .Y(n529) );
  INVX4 U776 ( .A(B[14]), .Y(n1059) );
  INVX1 U777 ( .A(n837), .Y(n838) );
  XNOR2X1 U778 ( .A(n530), .B(\SUMB[7][10] ), .Y(\SUMB[8][9] ) );
  XNOR2X1 U779 ( .A(\CARRYB[7][9] ), .B(\ab[8][9] ), .Y(n530) );
  NAND3X1 U780 ( .A(n665), .B(n663), .C(n664), .Y(n531) );
  INVX2 U781 ( .A(\SUMB[5][8] ), .Y(n742) );
  XNOR2X1 U782 ( .A(n318), .B(n532), .Y(n924) );
  NAND2X1 U783 ( .A(\SUMB[1][11] ), .B(n185), .Y(n533) );
  NAND2X1 U784 ( .A(\SUMB[1][11] ), .B(n104), .Y(n534) );
  NAND2X1 U785 ( .A(n104), .B(n185), .Y(n535) );
  NAND3X1 U786 ( .A(n535), .B(n533), .C(n534), .Y(\CARRYB[2][10] ) );
  INVX4 U787 ( .A(n1049), .Y(n579) );
  NAND3X1 U788 ( .A(n853), .B(n855), .C(n854), .Y(n536) );
  NAND3X1 U789 ( .A(n928), .B(n930), .C(n929), .Y(n537) );
  BUFX2 U790 ( .A(\SUMB[13][1] ), .Y(n538) );
  XNOR2X1 U791 ( .A(n539), .B(n82), .Y(\SUMB[4][11] ) );
  XNOR2X1 U792 ( .A(\CARRYB[3][11] ), .B(\ab[4][11] ), .Y(n539) );
  XOR2X1 U793 ( .A(n542), .B(n541), .Y(\SUMB[6][9] ) );
  INVX1 U794 ( .A(\SUMB[5][10] ), .Y(n542) );
  BUFX2 U795 ( .A(\CARRYB[12][0] ), .Y(n543) );
  BUFX2 U796 ( .A(\SUMB[7][2] ), .Y(n544) );
  NAND3X1 U797 ( .A(n923), .B(n922), .C(n921), .Y(n545) );
  NAND3X1 U798 ( .A(n850), .B(n851), .C(n852), .Y(n546) );
  XOR2X1 U799 ( .A(n547), .B(n137), .Y(\SUMB[15][1] ) );
  NAND2X1 U800 ( .A(\SUMB[14][2] ), .B(n321), .Y(n548) );
  NAND2X1 U801 ( .A(\SUMB[14][2] ), .B(\ab[15][1] ), .Y(n549) );
  NAND2X1 U802 ( .A(n321), .B(\ab[15][1] ), .Y(n550) );
  NAND3X1 U803 ( .A(n550), .B(n548), .C(n549), .Y(\CARRYB[15][1] ) );
  NAND2X1 U804 ( .A(\CARRYB[11][3] ), .B(\ab[12][3] ), .Y(n551) );
  NAND2X1 U805 ( .A(\SUMB[11][4] ), .B(\ab[12][3] ), .Y(n552) );
  NAND2X1 U806 ( .A(\SUMB[11][4] ), .B(\CARRYB[11][3] ), .Y(n553) );
  NAND3X1 U807 ( .A(n551), .B(n552), .C(n553), .Y(\CARRYB[12][3] ) );
  NAND2X1 U808 ( .A(\ab[13][2] ), .B(n324), .Y(n554) );
  NAND2X1 U809 ( .A(\SUMB[12][3] ), .B(\ab[13][2] ), .Y(n555) );
  NAND2X1 U810 ( .A(\SUMB[12][3] ), .B(n324), .Y(n556) );
  NAND3X1 U811 ( .A(n554), .B(n555), .C(n556), .Y(\CARRYB[13][2] ) );
  NAND2X1 U812 ( .A(n69), .B(\ab[2][9] ), .Y(n557) );
  NAND2X1 U813 ( .A(n69), .B(\SUMB[1][10] ), .Y(n558) );
  NAND2X1 U814 ( .A(\SUMB[1][10] ), .B(\ab[2][9] ), .Y(n559) );
  NAND3X1 U815 ( .A(n557), .B(n559), .C(n558), .Y(\CARRYB[2][9] ) );
  NAND2X1 U816 ( .A(\ab[3][8] ), .B(n396), .Y(n560) );
  NAND2X1 U817 ( .A(\SUMB[2][9] ), .B(\ab[3][8] ), .Y(n561) );
  NAND2X1 U818 ( .A(\SUMB[2][9] ), .B(n396), .Y(n562) );
  NAND3X1 U819 ( .A(n560), .B(n561), .C(n562), .Y(\CARRYB[3][8] ) );
  NAND2X1 U820 ( .A(n206), .B(n536), .Y(n563) );
  NAND2X1 U821 ( .A(\SUMB[7][6] ), .B(\ab[8][5] ), .Y(n564) );
  NAND2X1 U822 ( .A(n536), .B(\ab[8][5] ), .Y(n565) );
  NAND3X1 U823 ( .A(n565), .B(n563), .C(n564), .Y(\CARRYB[8][5] ) );
  NAND2X1 U824 ( .A(n943), .B(n945), .Y(n566) );
  NAND2X1 U825 ( .A(n944), .B(n567), .Y(n969) );
  INVX2 U826 ( .A(n566), .Y(n567) );
  XNOR2X1 U827 ( .A(n568), .B(n237), .Y(\SUMB[4][4] ) );
  XNOR2X1 U828 ( .A(\ab[4][4] ), .B(n266), .Y(n568) );
  XNOR2X1 U829 ( .A(n569), .B(n60), .Y(\SUMB[3][10] ) );
  XNOR2X1 U830 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .Y(n569) );
  XNOR2X1 U831 ( .A(n570), .B(\SUMB[13][5] ), .Y(\SUMB[14][4] ) );
  XNOR2X1 U832 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .Y(n570) );
  NAND3X1 U833 ( .A(n602), .B(n601), .C(n8), .Y(n571) );
  NAND2X1 U834 ( .A(n572), .B(n573), .Y(n574) );
  NAND2X1 U835 ( .A(n635), .B(n574), .Y(n578) );
  INVX1 U836 ( .A(\ab[5][2] ), .Y(n572) );
  XNOR2X1 U837 ( .A(n576), .B(n544), .Y(\SUMB[8][1] ) );
  XNOR2X1 U838 ( .A(\ab[8][1] ), .B(n428), .Y(n576) );
  XNOR2X1 U839 ( .A(n578), .B(n303), .Y(\SUMB[5][2] ) );
  INVX1 U840 ( .A(n1049), .Y(n1050) );
  INVX2 U841 ( .A(B[9]), .Y(n1049) );
  NAND3X1 U842 ( .A(n918), .B(n920), .C(n919), .Y(n580) );
  NAND3X1 U843 ( .A(n970), .B(n971), .C(n972), .Y(n581) );
  INVX4 U844 ( .A(n1063), .Y(n983) );
  NAND2X1 U845 ( .A(\SUMB[5][6] ), .B(n580), .Y(n582) );
  NAND2X1 U846 ( .A(\SUMB[5][6] ), .B(\ab[6][5] ), .Y(n583) );
  NAND2X1 U847 ( .A(n580), .B(\ab[6][5] ), .Y(n584) );
  NAND3X1 U848 ( .A(n583), .B(n584), .C(n582), .Y(\CARRYB[6][5] ) );
  NAND2X1 U849 ( .A(\ab[9][6] ), .B(n586), .Y(n587) );
  NAND2X1 U850 ( .A(\CARRYB[8][6] ), .B(n585), .Y(n588) );
  NAND2X1 U851 ( .A(n587), .B(n588), .Y(n956) );
  INVX1 U852 ( .A(\ab[9][6] ), .Y(n585) );
  INVX1 U853 ( .A(\CARRYB[8][6] ), .Y(n586) );
  NAND2X1 U854 ( .A(\SUMB[11][7] ), .B(\CARRYB[11][6] ), .Y(n591) );
  NAND2X1 U855 ( .A(\CARRYB[11][6] ), .B(\ab[12][6] ), .Y(n592) );
  NAND2X1 U856 ( .A(\SUMB[11][7] ), .B(\ab[12][6] ), .Y(n593) );
  NAND3X1 U857 ( .A(n592), .B(n591), .C(n593), .Y(\CARRYB[12][6] ) );
  NAND2X1 U858 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .Y(n595) );
  NAND2X1 U859 ( .A(\ab[4][4] ), .B(\SUMB[3][5] ), .Y(n596) );
  NAND2X1 U860 ( .A(\CARRYB[3][4] ), .B(\SUMB[3][5] ), .Y(n597) );
  NAND3X1 U861 ( .A(n595), .B(n596), .C(n597), .Y(\CARRYB[4][4] ) );
  NAND2X1 U862 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .Y(n598) );
  NAND2X1 U863 ( .A(\ab[5][3] ), .B(\SUMB[4][4] ), .Y(n599) );
  NAND2X1 U864 ( .A(\SUMB[4][4] ), .B(\CARRYB[4][3] ), .Y(n600) );
  NAND2X1 U865 ( .A(n419), .B(\SUMB[3][6] ), .Y(n601) );
  NAND2X1 U866 ( .A(\SUMB[3][6] ), .B(\ab[4][5] ), .Y(n602) );
  NAND2X1 U867 ( .A(n419), .B(\ab[4][5] ), .Y(n603) );
  NAND3X1 U868 ( .A(n602), .B(n603), .C(n601), .Y(\CARRYB[4][5] ) );
  XOR2X1 U869 ( .A(\SUMB[6][1] ), .B(\ab[7][0] ), .Y(n604) );
  XOR2X1 U870 ( .A(n661), .B(n604), .Y(\A1[5] ) );
  NAND2X1 U871 ( .A(n661), .B(\SUMB[6][1] ), .Y(n605) );
  NAND2X1 U872 ( .A(n661), .B(\ab[7][0] ), .Y(n606) );
  NAND2X1 U873 ( .A(\SUMB[6][1] ), .B(\ab[7][0] ), .Y(n607) );
  NAND3X1 U874 ( .A(n606), .B(n605), .C(n607), .Y(\CARRYB[7][0] ) );
  XOR2X1 U875 ( .A(\SUMB[3][2] ), .B(\ab[4][1] ), .Y(n608) );
  XOR2X1 U876 ( .A(\CARRYB[3][1] ), .B(n608), .Y(\SUMB[4][1] ) );
  NAND2X1 U877 ( .A(\CARRYB[3][1] ), .B(\SUMB[3][2] ), .Y(n609) );
  NAND2X1 U878 ( .A(\CARRYB[3][1] ), .B(\ab[4][1] ), .Y(n610) );
  NAND2X1 U879 ( .A(\SUMB[3][2] ), .B(\ab[4][1] ), .Y(n611) );
  NAND3X1 U880 ( .A(n610), .B(n609), .C(n611), .Y(\CARRYB[4][1] ) );
  XOR2X1 U881 ( .A(\ab[2][2] ), .B(n78), .Y(n612) );
  XOR2X1 U882 ( .A(n612), .B(\SUMB[1][3] ), .Y(\SUMB[2][2] ) );
  XOR2X1 U883 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .Y(n613) );
  XOR2X1 U884 ( .A(n613), .B(n205), .Y(\SUMB[3][1] ) );
  NAND2X1 U885 ( .A(\ab[2][2] ), .B(n78), .Y(n614) );
  NAND2X1 U886 ( .A(\ab[2][2] ), .B(\SUMB[1][3] ), .Y(n615) );
  NAND2X1 U887 ( .A(n78), .B(\SUMB[1][3] ), .Y(n616) );
  NAND3X1 U888 ( .A(n614), .B(n615), .C(n616), .Y(\CARRYB[2][2] ) );
  NAND2X1 U889 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .Y(n617) );
  NAND2X1 U890 ( .A(\ab[3][1] ), .B(\SUMB[2][2] ), .Y(n618) );
  NAND2X1 U891 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n619) );
  NAND3X1 U892 ( .A(n617), .B(n618), .C(n619), .Y(\CARRYB[3][1] ) );
  XOR2X1 U893 ( .A(\CARRYB[4][1] ), .B(\ab[5][1] ), .Y(n620) );
  XOR2X1 U894 ( .A(n625), .B(n620), .Y(\SUMB[5][1] ) );
  NAND2X1 U895 ( .A(\SUMB[4][2] ), .B(\CARRYB[4][1] ), .Y(n621) );
  NAND2X1 U896 ( .A(\SUMB[4][2] ), .B(\ab[5][1] ), .Y(n622) );
  NAND2X1 U897 ( .A(\CARRYB[4][1] ), .B(\ab[5][1] ), .Y(n623) );
  NAND3X1 U898 ( .A(n622), .B(n621), .C(n623), .Y(\CARRYB[5][1] ) );
  BUFX2 U899 ( .A(\SUMB[2][3] ), .Y(n624) );
  BUFX2 U900 ( .A(\SUMB[4][2] ), .Y(n625) );
  XNOR2X1 U901 ( .A(\CARRYB[6][6] ), .B(\ab[7][6] ), .Y(n626) );
  NAND2X1 U902 ( .A(\CARRYB[4][4] ), .B(\ab[5][4] ), .Y(n627) );
  NAND2X1 U903 ( .A(\SUMB[4][5] ), .B(\CARRYB[4][4] ), .Y(n628) );
  NAND2X1 U904 ( .A(\SUMB[4][5] ), .B(\ab[5][4] ), .Y(n629) );
  NAND3X1 U905 ( .A(n627), .B(n628), .C(n629), .Y(\CARRYB[5][4] ) );
  NAND2X1 U906 ( .A(\ab[6][3] ), .B(n56), .Y(n630) );
  NAND2X1 U907 ( .A(\SUMB[5][4] ), .B(\ab[6][3] ), .Y(n631) );
  NAND2X1 U908 ( .A(\SUMB[5][4] ), .B(n56), .Y(n632) );
  NAND3X1 U909 ( .A(n630), .B(n631), .C(n632), .Y(\CARRYB[6][3] ) );
  NAND3X1 U910 ( .A(n728), .B(n729), .C(n730), .Y(n633) );
  XOR2X1 U911 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .Y(n634) );
  XOR2X1 U912 ( .A(n634), .B(n17), .Y(\SUMB[6][1] ) );
  NAND2X1 U913 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .Y(n635) );
  NAND2X1 U914 ( .A(\ab[5][2] ), .B(\SUMB[4][3] ), .Y(n636) );
  NAND2X1 U915 ( .A(\SUMB[4][3] ), .B(\CARRYB[4][2] ), .Y(n637) );
  NAND3X1 U916 ( .A(n635), .B(n637), .C(n636), .Y(\CARRYB[5][2] ) );
  NAND2X1 U917 ( .A(\ab[6][1] ), .B(\SUMB[5][2] ), .Y(n638) );
  NAND2X1 U918 ( .A(\CARRYB[5][1] ), .B(\SUMB[5][2] ), .Y(n639) );
  NAND3X1 U919 ( .A(n203), .B(n638), .C(n639), .Y(\CARRYB[6][1] ) );
  INVX2 U920 ( .A(\ab[11][7] ), .Y(n654) );
  INVX2 U921 ( .A(\ab[4][7] ), .Y(n680) );
  NAND2X1 U922 ( .A(\SUMB[14][6] ), .B(\CARRYB[14][5] ), .Y(n640) );
  NAND2X1 U923 ( .A(\SUMB[14][6] ), .B(\ab[15][5] ), .Y(n641) );
  NAND2X1 U924 ( .A(\CARRYB[14][5] ), .B(\ab[15][5] ), .Y(n642) );
  NAND3X1 U925 ( .A(n641), .B(n640), .C(n642), .Y(\CARRYB[15][5] ) );
  XOR2X1 U926 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .Y(n643) );
  XOR2X1 U927 ( .A(n643), .B(\SUMB[13][7] ), .Y(\SUMB[14][6] ) );
  NAND2X1 U928 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .Y(n644) );
  NAND2X1 U929 ( .A(\ab[13][7] ), .B(\SUMB[12][8] ), .Y(n645) );
  NAND2X1 U930 ( .A(\CARRYB[12][7] ), .B(\SUMB[12][8] ), .Y(n646) );
  NAND3X1 U931 ( .A(n644), .B(n646), .C(n645), .Y(\CARRYB[13][7] ) );
  NAND2X1 U932 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .Y(n647) );
  NAND2X1 U933 ( .A(\SUMB[13][7] ), .B(\ab[14][6] ), .Y(n648) );
  NAND2X1 U934 ( .A(\SUMB[13][7] ), .B(\CARRYB[13][6] ), .Y(n649) );
  NAND3X1 U935 ( .A(n647), .B(n648), .C(n649), .Y(\CARRYB[14][6] ) );
  XOR2X1 U936 ( .A(\CARRYB[11][7] ), .B(\ab[12][7] ), .Y(n650) );
  XOR2X1 U937 ( .A(\SUMB[11][8] ), .B(n650), .Y(\SUMB[12][7] ) );
  NAND2X1 U938 ( .A(\SUMB[11][8] ), .B(n229), .Y(n651) );
  NAND2X1 U939 ( .A(\SUMB[11][8] ), .B(\ab[12][7] ), .Y(n652) );
  NAND2X1 U940 ( .A(n229), .B(\ab[12][7] ), .Y(n653) );
  NAND3X1 U941 ( .A(n652), .B(n651), .C(n653), .Y(\CARRYB[12][7] ) );
  INVX1 U942 ( .A(n1043), .Y(n1089) );
  INVX1 U943 ( .A(n657), .Y(n658) );
  INVX4 U944 ( .A(B[5]), .Y(n1042) );
  BUFX2 U945 ( .A(\CARRYB[3][7] ), .Y(n655) );
  NAND3X1 U946 ( .A(n940), .B(n941), .C(n942), .Y(n656) );
  INVX2 U947 ( .A(\SUMB[7][3] ), .Y(n674) );
  NAND3X1 U948 ( .A(n423), .B(n1009), .C(n1010), .Y(n659) );
  INVX4 U949 ( .A(B[6]), .Y(n1044) );
  OR2X2 U950 ( .A(n464), .B(n1028), .Y(n703) );
  BUFX4 U951 ( .A(\CARRYB[6][0] ), .Y(n661) );
  INVX4 U952 ( .A(B[3]), .Y(n1038) );
  XOR2X1 U953 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U954 ( .A(\CARRYB[3][3] ), .B(\ab[4][3] ), .Y(n662) );
  XOR2X1 U955 ( .A(n438), .B(n662), .Y(\SUMB[4][3] ) );
  NAND2X1 U956 ( .A(\SUMB[3][4] ), .B(n145), .Y(n663) );
  NAND2X1 U957 ( .A(\SUMB[3][4] ), .B(\ab[4][3] ), .Y(n664) );
  NAND2X1 U958 ( .A(n145), .B(\ab[4][3] ), .Y(n665) );
  NAND3X1 U959 ( .A(n664), .B(n663), .C(n665), .Y(\CARRYB[4][3] ) );
  XOR2X1 U960 ( .A(n144), .B(\ab[6][2] ), .Y(n667) );
  XOR2X1 U961 ( .A(n417), .B(n667), .Y(\SUMB[6][2] ) );
  NAND2X1 U962 ( .A(\CARRYB[5][2] ), .B(\SUMB[5][3] ), .Y(n668) );
  NAND2X1 U963 ( .A(\SUMB[5][3] ), .B(\ab[6][2] ), .Y(n669) );
  NAND2X1 U964 ( .A(\CARRYB[5][2] ), .B(\ab[6][2] ), .Y(n670) );
  NAND3X1 U965 ( .A(n670), .B(n669), .C(n668), .Y(\CARRYB[6][2] ) );
  NAND2X1 U966 ( .A(n675), .B(\CARRYB[6][2] ), .Y(n671) );
  NAND2X1 U967 ( .A(\ab[7][2] ), .B(n1027), .Y(n672) );
  NAND2X1 U968 ( .A(n671), .B(n672), .Y(n1008) );
  INVX1 U969 ( .A(\ab[7][2] ), .Y(n675) );
  XOR2X1 U970 ( .A(n673), .B(n674), .Y(\SUMB[8][2] ) );
  INVX4 U971 ( .A(B[0]), .Y(n1032) );
  INVX1 U972 ( .A(\SUMB[6][4] ), .Y(n676) );
  XNOR2X1 U973 ( .A(n633), .B(\ab[9][2] ), .Y(n677) );
  NAND3X1 U974 ( .A(n783), .B(n784), .C(n785), .Y(n678) );
  NAND3X1 U975 ( .A(n842), .B(n841), .C(n843), .Y(n679) );
  XOR2X1 U976 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .Y(n681) );
  XOR2X1 U977 ( .A(n681), .B(n162), .Y(\SUMB[4][12] ) );
  NAND2X1 U978 ( .A(\ab[4][12] ), .B(n128), .Y(n682) );
  NAND2X1 U979 ( .A(\ab[4][12] ), .B(\SUMB[3][13] ), .Y(n683) );
  NAND2X1 U980 ( .A(n128), .B(\SUMB[3][13] ), .Y(n684) );
  NAND3X1 U981 ( .A(n682), .B(n683), .C(n684), .Y(\CARRYB[4][12] ) );
  NAND2X1 U982 ( .A(\ab[5][11] ), .B(n832), .Y(n685) );
  NAND2X1 U983 ( .A(\ab[5][11] ), .B(\SUMB[4][12] ), .Y(n686) );
  NAND2X1 U984 ( .A(n832), .B(\SUMB[4][12] ), .Y(n687) );
  NAND3X1 U985 ( .A(n685), .B(n686), .C(n687), .Y(\CARRYB[5][11] ) );
  NAND2X1 U986 ( .A(\ab[14][7] ), .B(n221), .Y(n688) );
  NAND2X1 U987 ( .A(\ab[14][7] ), .B(\SUMB[13][8] ), .Y(n689) );
  NAND2X1 U988 ( .A(n221), .B(\SUMB[13][8] ), .Y(n690) );
  NAND3X1 U989 ( .A(n688), .B(n689), .C(n690), .Y(\CARRYB[14][7] ) );
  NAND2X1 U990 ( .A(\ab[15][6] ), .B(n269), .Y(n691) );
  NAND2X1 U991 ( .A(\ab[15][6] ), .B(\SUMB[14][7] ), .Y(n692) );
  NAND2X1 U992 ( .A(n269), .B(\SUMB[14][7] ), .Y(n693) );
  NAND3X1 U993 ( .A(n691), .B(n692), .C(n693), .Y(\CARRYB[15][6] ) );
  NAND2X1 U994 ( .A(\ab[11][9] ), .B(n135), .Y(n694) );
  NAND2X1 U995 ( .A(\ab[11][9] ), .B(\SUMB[10][10] ), .Y(n695) );
  NAND2X1 U996 ( .A(n135), .B(\SUMB[10][10] ), .Y(n696) );
  NAND3X1 U997 ( .A(n694), .B(n695), .C(n696), .Y(\CARRYB[11][9] ) );
  XOR2X1 U998 ( .A(\ab[12][9] ), .B(\SUMB[11][10] ), .Y(n697) );
  XOR2X1 U999 ( .A(n697), .B(\CARRYB[11][9] ), .Y(\SUMB[12][9] ) );
  NAND2X1 U1000 ( .A(\ab[12][9] ), .B(\SUMB[11][10] ), .Y(n698) );
  NAND2X1 U1001 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .Y(n699) );
  NAND2X1 U1002 ( .A(\SUMB[11][10] ), .B(\CARRYB[11][9] ), .Y(n700) );
  NAND3X1 U1003 ( .A(n698), .B(n699), .C(n700), .Y(\CARRYB[12][9] ) );
  INVX2 U1004 ( .A(\CARRYB[2][4] ), .Y(n701) );
  XOR2X1 U1005 ( .A(n702), .B(\SUMB[11][3] ), .Y(\SUMB[12][2] ) );
  NAND2X1 U1006 ( .A(\SUMB[10][4] ), .B(\ab[11][3] ), .Y(n704) );
  NAND2X1 U1007 ( .A(n1029), .B(\SUMB[10][4] ), .Y(n705) );
  NAND3X1 U1008 ( .A(n703), .B(n705), .C(n704), .Y(\CARRYB[11][3] ) );
  NAND2X1 U1009 ( .A(n316), .B(\ab[12][2] ), .Y(n706) );
  NAND2X1 U1010 ( .A(\SUMB[11][3] ), .B(\ab[12][2] ), .Y(n707) );
  NAND2X1 U1011 ( .A(n316), .B(\SUMB[11][3] ), .Y(n708) );
  NAND3X1 U1012 ( .A(n706), .B(n707), .C(n708), .Y(\CARRYB[12][2] ) );
  NAND2X1 U1013 ( .A(\ab[3][9] ), .B(n341), .Y(n709) );
  NAND2X1 U1014 ( .A(\SUMB[2][10] ), .B(\ab[3][9] ), .Y(n710) );
  NAND2X1 U1015 ( .A(\SUMB[2][10] ), .B(n341), .Y(n711) );
  NAND3X1 U1016 ( .A(n709), .B(n710), .C(n711), .Y(\CARRYB[3][9] ) );
  NAND2X1 U1017 ( .A(n914), .B(\ab[4][8] ), .Y(n712) );
  NAND2X1 U1018 ( .A(\SUMB[3][9] ), .B(\ab[4][8] ), .Y(n713) );
  NAND2X1 U1019 ( .A(\SUMB[3][9] ), .B(n914), .Y(n714) );
  NAND3X1 U1020 ( .A(n712), .B(n713), .C(n714), .Y(\CARRYB[4][8] ) );
  XOR2X1 U1021 ( .A(n715), .B(n742), .Y(\SUMB[6][7] ) );
  INVX1 U1022 ( .A(n1052), .Y(n1085) );
  INVX2 U1023 ( .A(\SUMB[1][9] ), .Y(n722) );
  NAND2X1 U1024 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .Y(n716) );
  NAND2X1 U1025 ( .A(\SUMB[8][3] ), .B(\ab[9][2] ), .Y(n717) );
  NAND2X1 U1026 ( .A(\CARRYB[8][2] ), .B(\SUMB[8][3] ), .Y(n718) );
  NAND3X1 U1027 ( .A(n716), .B(n717), .C(n718), .Y(\CARRYB[9][2] ) );
  NAND2X1 U1028 ( .A(\ab[10][1] ), .B(n1026), .Y(n719) );
  NAND2X1 U1029 ( .A(\ab[10][1] ), .B(\SUMB[9][2] ), .Y(n720) );
  NAND2X1 U1030 ( .A(n1026), .B(\SUMB[9][2] ), .Y(n721) );
  NAND3X1 U1031 ( .A(n719), .B(n720), .C(n721), .Y(\CARRYB[10][1] ) );
  NAND3X1 U1032 ( .A(n975), .B(n974), .C(n18), .Y(n723) );
  NAND2X1 U1033 ( .A(n436), .B(\ab[7][3] ), .Y(n725) );
  NAND2X1 U1034 ( .A(\SUMB[6][4] ), .B(n436), .Y(n726) );
  NAND2X1 U1035 ( .A(\SUMB[6][4] ), .B(\ab[7][3] ), .Y(n727) );
  NAND3X1 U1036 ( .A(n725), .B(n727), .C(n726), .Y(\CARRYB[7][3] ) );
  NAND2X1 U1037 ( .A(\ab[8][2] ), .B(n659), .Y(n728) );
  NAND2X1 U1038 ( .A(\SUMB[7][3] ), .B(\ab[8][2] ), .Y(n729) );
  NAND2X1 U1039 ( .A(n659), .B(\SUMB[7][3] ), .Y(n730) );
  NAND3X1 U1040 ( .A(n728), .B(n729), .C(n730), .Y(\CARRYB[8][2] ) );
  INVX1 U1041 ( .A(n1047), .Y(n1087) );
  XOR2X1 U1042 ( .A(\SUMB[1][4] ), .B(\ab[2][3] ), .Y(n732) );
  XOR2X1 U1043 ( .A(n732), .B(n1021), .Y(\SUMB[2][3] ) );
  NAND2X1 U1044 ( .A(\SUMB[1][4] ), .B(n1021), .Y(n733) );
  NAND2X1 U1045 ( .A(n1021), .B(\ab[2][3] ), .Y(n734) );
  NAND2X1 U1046 ( .A(\SUMB[1][4] ), .B(\ab[2][3] ), .Y(n735) );
  NAND3X1 U1047 ( .A(n734), .B(n733), .C(n735), .Y(\CARRYB[2][3] ) );
  INVX4 U1048 ( .A(A[2]), .Y(n1064) );
  NOR2X1 U1049 ( .A(n1061), .B(n1044), .Y(\ab[0][6] ) );
  NAND2X1 U1050 ( .A(n263), .B(\ab[10][5] ), .Y(n736) );
  NAND2X1 U1051 ( .A(\SUMB[9][6] ), .B(\ab[10][5] ), .Y(n737) );
  NAND2X1 U1052 ( .A(\SUMB[9][6] ), .B(n263), .Y(n738) );
  NAND3X1 U1053 ( .A(n736), .B(n737), .C(n738), .Y(\CARRYB[10][5] ) );
  NAND2X1 U1054 ( .A(n395), .B(\ab[11][4] ), .Y(n739) );
  NAND2X1 U1055 ( .A(\SUMB[10][5] ), .B(\ab[11][4] ), .Y(n740) );
  NAND2X1 U1056 ( .A(n395), .B(\SUMB[10][5] ), .Y(n741) );
  NAND3X1 U1057 ( .A(n739), .B(n740), .C(n741), .Y(\CARRYB[11][4] ) );
  NAND2X1 U1058 ( .A(n340), .B(\ab[12][4] ), .Y(n743) );
  NAND2X1 U1059 ( .A(\ab[12][4] ), .B(\SUMB[11][5] ), .Y(n744) );
  NAND2X1 U1060 ( .A(n340), .B(\SUMB[11][5] ), .Y(n745) );
  NAND3X1 U1061 ( .A(n743), .B(n744), .C(n745), .Y(\CARRYB[12][4] ) );
  NAND2X1 U1062 ( .A(\SUMB[12][5] ), .B(\ab[13][4] ), .Y(n746) );
  NAND2X1 U1063 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .Y(n747) );
  NAND2X1 U1064 ( .A(\SUMB[12][5] ), .B(\CARRYB[12][4] ), .Y(n748) );
  NAND3X1 U1065 ( .A(n746), .B(n747), .C(n748), .Y(\CARRYB[13][4] ) );
  INVX1 U1066 ( .A(n579), .Y(n1086) );
  XNOR2X1 U1067 ( .A(\SUMB[15][1] ), .B(n749), .Y(\A1[14] ) );
  NOR2X1 U1068 ( .A(n1061), .B(n1048), .Y(\ab[0][8] ) );
  NAND2X1 U1069 ( .A(\SUMB[13][4] ), .B(\CARRYB[13][3] ), .Y(n750) );
  NAND2X1 U1070 ( .A(\SUMB[13][4] ), .B(\ab[14][3] ), .Y(n751) );
  NAND2X1 U1071 ( .A(n678), .B(\ab[14][3] ), .Y(n752) );
  NAND3X1 U1072 ( .A(n752), .B(n751), .C(n750), .Y(\CARRYB[14][3] ) );
  NAND2X1 U1073 ( .A(\ab[3][10] ), .B(n134), .Y(n753) );
  NAND2X1 U1074 ( .A(\SUMB[2][11] ), .B(\ab[3][10] ), .Y(n754) );
  NAND2X1 U1075 ( .A(\SUMB[2][11] ), .B(n134), .Y(n755) );
  NAND3X1 U1076 ( .A(n753), .B(n754), .C(n755), .Y(\CARRYB[3][10] ) );
  NAND2X1 U1077 ( .A(\ab[4][9] ), .B(n389), .Y(n756) );
  NAND2X1 U1078 ( .A(\SUMB[3][10] ), .B(\ab[4][9] ), .Y(n757) );
  NAND2X1 U1079 ( .A(\SUMB[3][10] ), .B(n389), .Y(n758) );
  NAND3X1 U1080 ( .A(n756), .B(n757), .C(n758), .Y(\CARRYB[4][9] ) );
  NAND2X1 U1081 ( .A(\ab[11][6] ), .B(n307), .Y(n759) );
  NAND2X1 U1082 ( .A(\SUMB[10][7] ), .B(\ab[11][6] ), .Y(n760) );
  NAND2X1 U1083 ( .A(\SUMB[10][7] ), .B(n307), .Y(n761) );
  NAND3X1 U1084 ( .A(n759), .B(n760), .C(n761), .Y(\CARRYB[11][6] ) );
  NAND2X1 U1085 ( .A(\ab[12][5] ), .B(n232), .Y(n762) );
  NAND2X1 U1086 ( .A(\SUMB[11][6] ), .B(\ab[12][5] ), .Y(n763) );
  NAND2X1 U1087 ( .A(\SUMB[11][6] ), .B(n232), .Y(n764) );
  NAND3X1 U1088 ( .A(n762), .B(n763), .C(n764), .Y(\CARRYB[12][5] ) );
  XOR2X1 U1089 ( .A(\CARRYB[7][11] ), .B(\ab[8][11] ), .Y(n765) );
  XOR2X1 U1090 ( .A(n765), .B(\SUMB[7][12] ), .Y(\SUMB[8][11] ) );
  NAND2X1 U1091 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .Y(n766) );
  NAND2X1 U1092 ( .A(\ab[8][11] ), .B(\SUMB[7][12] ), .Y(n767) );
  NAND2X1 U1093 ( .A(\CARRYB[7][11] ), .B(\SUMB[7][12] ), .Y(n768) );
  NAND3X1 U1094 ( .A(n766), .B(n767), .C(n768), .Y(\CARRYB[8][11] ) );
  NAND2X1 U1095 ( .A(\ab[9][10] ), .B(n111), .Y(n769) );
  NAND2X1 U1096 ( .A(\ab[9][10] ), .B(\SUMB[8][11] ), .Y(n770) );
  NAND2X1 U1097 ( .A(n111), .B(\SUMB[8][11] ), .Y(n771) );
  NAND3X1 U1098 ( .A(n769), .B(n770), .C(n771), .Y(\CARRYB[9][10] ) );
  XOR2X1 U1099 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .Y(n772) );
  XOR2X1 U1100 ( .A(n772), .B(\SUMB[12][7] ), .Y(\SUMB[13][6] ) );
  NAND2X1 U1101 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .Y(n773) );
  NAND2X1 U1102 ( .A(\SUMB[12][7] ), .B(\ab[13][6] ), .Y(n774) );
  NAND2X1 U1103 ( .A(\CARRYB[12][6] ), .B(\SUMB[12][7] ), .Y(n775) );
  NAND3X1 U1104 ( .A(n773), .B(n774), .C(n775), .Y(\CARRYB[13][6] ) );
  NAND2X1 U1105 ( .A(\ab[14][5] ), .B(n326), .Y(n776) );
  NAND2X1 U1106 ( .A(\SUMB[13][6] ), .B(\ab[14][5] ), .Y(n777) );
  NAND2X1 U1107 ( .A(n326), .B(\SUMB[13][6] ), .Y(n778) );
  NAND3X1 U1108 ( .A(n776), .B(n777), .C(n778), .Y(\CARRYB[14][5] ) );
  XOR2X1 U1109 ( .A(n779), .B(\SUMB[1][14] ), .Y(\SUMB[2][13] ) );
  NAND2X1 U1110 ( .A(\SUMB[1][14] ), .B(\CARRYB[1][13] ), .Y(n780) );
  NAND2X1 U1111 ( .A(\SUMB[1][14] ), .B(\ab[2][13] ), .Y(n781) );
  NAND2X1 U1112 ( .A(\CARRYB[1][13] ), .B(\ab[2][13] ), .Y(n782) );
  NAND3X1 U1113 ( .A(n782), .B(n780), .C(n781), .Y(\CARRYB[2][13] ) );
  NAND2X1 U1114 ( .A(\SUMB[12][4] ), .B(\ab[13][3] ), .Y(n784) );
  NAND2X1 U1115 ( .A(\SUMB[12][4] ), .B(n798), .Y(n785) );
  NAND3X1 U1116 ( .A(n783), .B(n784), .C(n785), .Y(\CARRYB[13][3] ) );
  NAND2X1 U1117 ( .A(\CARRYB[13][2] ), .B(\ab[14][2] ), .Y(n786) );
  NAND2X1 U1118 ( .A(\SUMB[13][3] ), .B(\ab[14][2] ), .Y(n787) );
  NAND2X1 U1119 ( .A(\SUMB[13][3] ), .B(\CARRYB[13][2] ), .Y(n788) );
  NAND3X1 U1120 ( .A(n786), .B(n787), .C(n788), .Y(\CARRYB[14][2] ) );
  NAND2X1 U1121 ( .A(\SUMB[4][9] ), .B(n451), .Y(n789) );
  NAND2X1 U1122 ( .A(\SUMB[4][9] ), .B(\ab[5][8] ), .Y(n790) );
  NAND2X1 U1123 ( .A(n451), .B(\ab[5][8] ), .Y(n791) );
  NAND3X1 U1124 ( .A(n791), .B(n789), .C(n790), .Y(\CARRYB[5][8] ) );
  NAND3X1 U1125 ( .A(n901), .B(n903), .C(n902), .Y(n792) );
  XOR2X1 U1126 ( .A(n32), .B(\ab[13][0] ), .Y(n793) );
  XOR2X1 U1127 ( .A(n543), .B(n793), .Y(\A1[11] ) );
  NAND2X1 U1128 ( .A(\SUMB[12][1] ), .B(\CARRYB[12][0] ), .Y(n794) );
  NAND2X1 U1129 ( .A(\CARRYB[12][0] ), .B(\ab[13][0] ), .Y(n795) );
  NAND2X1 U1130 ( .A(\SUMB[12][1] ), .B(\ab[13][0] ), .Y(n796) );
  NAND3X1 U1131 ( .A(n795), .B(n796), .C(n794), .Y(\CARRYB[13][0] ) );
  INVX2 U1132 ( .A(\CARRYB[12][3] ), .Y(n797) );
  NAND2X1 U1133 ( .A(\ab[6][9] ), .B(n836), .Y(n799) );
  NAND2X1 U1134 ( .A(\SUMB[5][10] ), .B(\ab[6][9] ), .Y(n800) );
  NAND2X1 U1135 ( .A(\SUMB[5][10] ), .B(n836), .Y(n801) );
  NAND3X1 U1136 ( .A(n800), .B(n799), .C(n801), .Y(\CARRYB[6][9] ) );
  NAND2X1 U1137 ( .A(\ab[7][8] ), .B(n656), .Y(n802) );
  NAND2X1 U1138 ( .A(\ab[7][8] ), .B(\SUMB[6][9] ), .Y(n803) );
  NAND2X1 U1139 ( .A(n656), .B(\SUMB[6][9] ), .Y(n804) );
  NAND3X1 U1140 ( .A(n802), .B(n803), .C(n804), .Y(\CARRYB[7][8] ) );
  NAND2X1 U1141 ( .A(\ab[6][10] ), .B(n838), .Y(n805) );
  NAND2X1 U1142 ( .A(\ab[6][10] ), .B(\SUMB[5][11] ), .Y(n806) );
  NAND2X1 U1143 ( .A(n838), .B(\SUMB[5][11] ), .Y(n807) );
  NAND3X1 U1144 ( .A(n805), .B(n806), .C(n807), .Y(\CARRYB[6][10] ) );
  NAND2X1 U1145 ( .A(\ab[7][9] ), .B(n840), .Y(n808) );
  NAND2X1 U1146 ( .A(\ab[7][9] ), .B(\SUMB[6][10] ), .Y(n809) );
  NAND2X1 U1147 ( .A(n840), .B(\SUMB[6][10] ), .Y(n810) );
  NAND3X1 U1148 ( .A(n808), .B(n809), .C(n810), .Y(\CARRYB[7][9] ) );
  NAND2X1 U1149 ( .A(\ab[3][11] ), .B(n184), .Y(n811) );
  NAND2X1 U1150 ( .A(\SUMB[2][12] ), .B(\ab[3][11] ), .Y(n812) );
  NAND2X1 U1151 ( .A(\SUMB[2][12] ), .B(n184), .Y(n813) );
  NAND3X1 U1152 ( .A(n811), .B(n812), .C(n813), .Y(\CARRYB[3][11] ) );
  NAND2X1 U1153 ( .A(\ab[4][10] ), .B(n834), .Y(n814) );
  NAND2X1 U1154 ( .A(\SUMB[3][11] ), .B(\ab[4][10] ), .Y(n815) );
  NAND2X1 U1155 ( .A(\SUMB[3][11] ), .B(n834), .Y(n816) );
  NAND3X1 U1156 ( .A(n814), .B(n815), .C(n816), .Y(\CARRYB[4][10] ) );
  NAND2X1 U1157 ( .A(\ab[7][10] ), .B(n313), .Y(n817) );
  NAND2X1 U1158 ( .A(\ab[7][10] ), .B(\SUMB[6][11] ), .Y(n818) );
  NAND2X1 U1159 ( .A(n313), .B(\SUMB[6][11] ), .Y(n819) );
  NAND3X1 U1160 ( .A(n817), .B(n818), .C(n819), .Y(\CARRYB[7][10] ) );
  NAND2X1 U1161 ( .A(\ab[8][9] ), .B(n327), .Y(n820) );
  NAND2X1 U1162 ( .A(\ab[8][9] ), .B(\SUMB[7][10] ), .Y(n821) );
  NAND2X1 U1163 ( .A(n327), .B(\SUMB[7][10] ), .Y(n822) );
  NAND3X1 U1164 ( .A(n820), .B(n821), .C(n822), .Y(\CARRYB[8][9] ) );
  NAND2X1 U1165 ( .A(\ab[3][12] ), .B(n116), .Y(n823) );
  NAND2X1 U1166 ( .A(\SUMB[2][13] ), .B(\ab[3][12] ), .Y(n824) );
  NAND2X1 U1167 ( .A(\SUMB[2][13] ), .B(n116), .Y(n825) );
  NAND3X1 U1168 ( .A(n823), .B(n824), .C(n825), .Y(\CARRYB[3][12] ) );
  NAND2X1 U1169 ( .A(\ab[4][11] ), .B(n268), .Y(n826) );
  NAND2X1 U1170 ( .A(\SUMB[3][12] ), .B(\ab[4][11] ), .Y(n827) );
  NAND2X1 U1171 ( .A(\SUMB[3][12] ), .B(n268), .Y(n828) );
  NAND3X1 U1172 ( .A(n826), .B(n827), .C(n828), .Y(\CARRYB[4][11] ) );
  INVX2 U1173 ( .A(\CARRYB[4][12] ), .Y(n829) );
  INVX2 U1174 ( .A(\CARRYB[4][11] ), .Y(n831) );
  INVX2 U1175 ( .A(\CARRYB[5][9] ), .Y(n835) );
  INVX2 U1176 ( .A(\CARRYB[5][10] ), .Y(n837) );
  NAND2X1 U1177 ( .A(n165), .B(\ab[5][7] ), .Y(n841) );
  NAND2X1 U1178 ( .A(\SUMB[4][8] ), .B(\ab[5][7] ), .Y(n842) );
  NAND2X1 U1179 ( .A(\SUMB[4][8] ), .B(n165), .Y(n843) );
  NAND3X1 U1180 ( .A(n842), .B(n841), .C(n843), .Y(\CARRYB[5][7] ) );
  NAND2X1 U1181 ( .A(\ab[6][6] ), .B(n537), .Y(n844) );
  NAND2X1 U1182 ( .A(\SUMB[5][7] ), .B(\ab[6][6] ), .Y(n845) );
  NAND2X1 U1183 ( .A(n537), .B(\SUMB[5][7] ), .Y(n846) );
  NAND3X1 U1184 ( .A(n844), .B(n845), .C(n846), .Y(\CARRYB[6][6] ) );
  NAND2X1 U1185 ( .A(n442), .B(\ab[11][2] ), .Y(n847) );
  NAND2X1 U1186 ( .A(\ab[11][2] ), .B(\SUMB[10][3] ), .Y(n848) );
  NAND2X1 U1187 ( .A(n442), .B(\SUMB[10][3] ), .Y(n849) );
  NAND3X1 U1188 ( .A(n847), .B(n848), .C(n849), .Y(\CARRYB[11][2] ) );
  NAND2X1 U1189 ( .A(n594), .B(\ab[12][1] ), .Y(n850) );
  NAND2X1 U1190 ( .A(\SUMB[11][2] ), .B(\ab[12][1] ), .Y(n851) );
  NAND2X1 U1191 ( .A(\SUMB[11][2] ), .B(n594), .Y(n852) );
  NAND3X1 U1192 ( .A(n851), .B(n850), .C(n852), .Y(\CARRYB[12][1] ) );
  NAND2X1 U1193 ( .A(\ab[7][5] ), .B(n323), .Y(n853) );
  NAND2X1 U1194 ( .A(\SUMB[6][6] ), .B(\ab[7][5] ), .Y(n854) );
  NAND2X1 U1195 ( .A(\SUMB[6][6] ), .B(n323), .Y(n855) );
  NAND3X1 U1196 ( .A(n853), .B(n854), .C(n855), .Y(\CARRYB[7][5] ) );
  NAND2X1 U1197 ( .A(\ab[8][4] ), .B(n581), .Y(n856) );
  NAND2X1 U1198 ( .A(\SUMB[7][5] ), .B(\ab[8][4] ), .Y(n857) );
  NAND2X1 U1199 ( .A(\SUMB[7][5] ), .B(n581), .Y(n858) );
  NAND3X1 U1200 ( .A(n856), .B(n857), .C(n858), .Y(\CARRYB[8][4] ) );
  XOR2X1 U1201 ( .A(n265), .B(\ab[14][0] ), .Y(n859) );
  XOR2X1 U1202 ( .A(n859), .B(n538), .Y(\A1[12] ) );
  NAND2X1 U1203 ( .A(n546), .B(\ab[13][1] ), .Y(n860) );
  NAND2X1 U1204 ( .A(\SUMB[12][2] ), .B(\ab[13][1] ), .Y(n861) );
  NAND2X1 U1205 ( .A(\SUMB[12][2] ), .B(n546), .Y(n862) );
  NAND3X1 U1206 ( .A(n860), .B(n861), .C(n862), .Y(\CARRYB[13][1] ) );
  NAND2X1 U1207 ( .A(\CARRYB[13][0] ), .B(\ab[14][0] ), .Y(n863) );
  NAND2X1 U1208 ( .A(\SUMB[13][1] ), .B(\ab[14][0] ), .Y(n864) );
  NAND2X1 U1209 ( .A(\SUMB[13][1] ), .B(\CARRYB[13][0] ), .Y(n865) );
  NAND3X1 U1210 ( .A(n864), .B(n865), .C(n863), .Y(\CARRYB[14][0] ) );
  NAND2X1 U1211 ( .A(\ab[9][7] ), .B(n494), .Y(n868) );
  NAND2X1 U1212 ( .A(\SUMB[8][8] ), .B(\ab[9][7] ), .Y(n869) );
  NAND2X1 U1213 ( .A(\SUMB[8][8] ), .B(n494), .Y(n870) );
  NAND3X1 U1214 ( .A(n868), .B(n869), .C(n870), .Y(\CARRYB[9][7] ) );
  NAND2X1 U1215 ( .A(\ab[10][6] ), .B(n422), .Y(n871) );
  NAND2X1 U1216 ( .A(\SUMB[9][7] ), .B(\ab[10][6] ), .Y(n872) );
  NAND2X1 U1217 ( .A(\SUMB[9][7] ), .B(n422), .Y(n873) );
  NAND3X1 U1218 ( .A(n871), .B(n872), .C(n873), .Y(\CARRYB[10][6] ) );
  XOR2X1 U1219 ( .A(n874), .B(n43), .Y(\SUMB[3][13] ) );
  NAND2X1 U1220 ( .A(\ab[2][14] ), .B(n195), .Y(n875) );
  NAND2X1 U1221 ( .A(\ab[2][14] ), .B(\ab[1][15] ), .Y(n876) );
  NAND2X1 U1222 ( .A(n195), .B(\ab[1][15] ), .Y(n877) );
  NAND3X1 U1223 ( .A(n875), .B(n876), .C(n877), .Y(\CARRYB[2][14] ) );
  NAND2X1 U1224 ( .A(\ab[3][13] ), .B(n163), .Y(n878) );
  NAND2X1 U1225 ( .A(\ab[3][13] ), .B(\SUMB[2][14] ), .Y(n879) );
  NAND2X1 U1226 ( .A(n163), .B(\SUMB[2][14] ), .Y(n880) );
  NAND3X1 U1227 ( .A(n878), .B(n879), .C(n880), .Y(\CARRYB[3][13] ) );
  NAND2X1 U1228 ( .A(\ab[10][8] ), .B(n328), .Y(n881) );
  NAND2X1 U1229 ( .A(\SUMB[9][9] ), .B(\ab[10][8] ), .Y(n882) );
  NAND2X1 U1230 ( .A(n328), .B(\SUMB[9][9] ), .Y(n883) );
  NAND3X1 U1231 ( .A(n881), .B(n882), .C(n883), .Y(\CARRYB[10][8] ) );
  NAND2X1 U1232 ( .A(\ab[11][7] ), .B(n658), .Y(n884) );
  NAND2X1 U1233 ( .A(\SUMB[10][8] ), .B(\ab[11][7] ), .Y(n885) );
  NAND2X1 U1234 ( .A(\SUMB[10][8] ), .B(n658), .Y(n886) );
  NAND3X1 U1235 ( .A(n884), .B(n885), .C(n886), .Y(\CARRYB[11][7] ) );
  XOR2X1 U1236 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .Y(n887) );
  XOR2X1 U1237 ( .A(n887), .B(\SUMB[12][6] ), .Y(\SUMB[13][5] ) );
  NAND2X1 U1238 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .Y(n888) );
  NAND2X1 U1239 ( .A(\SUMB[12][6] ), .B(\ab[13][5] ), .Y(n889) );
  NAND2X1 U1240 ( .A(\SUMB[12][6] ), .B(\CARRYB[12][5] ), .Y(n890) );
  NAND3X1 U1241 ( .A(n888), .B(n889), .C(n890), .Y(\CARRYB[13][5] ) );
  NAND2X1 U1242 ( .A(\ab[14][4] ), .B(n495), .Y(n891) );
  NAND2X1 U1243 ( .A(\SUMB[13][5] ), .B(\ab[14][4] ), .Y(n892) );
  NAND2X1 U1244 ( .A(n495), .B(\SUMB[13][5] ), .Y(n893) );
  NAND3X1 U1245 ( .A(n891), .B(n892), .C(n893), .Y(\CARRYB[14][4] ) );
  INVX1 U1246 ( .A(n1061), .Y(n894) );
  NAND2X1 U1247 ( .A(\ab[9][5] ), .B(n393), .Y(n895) );
  NAND2X1 U1248 ( .A(\SUMB[8][6] ), .B(\ab[9][5] ), .Y(n896) );
  NAND2X1 U1249 ( .A(n393), .B(\SUMB[8][6] ), .Y(n897) );
  NAND3X1 U1250 ( .A(n895), .B(n896), .C(n897), .Y(\CARRYB[9][5] ) );
  NAND2X1 U1251 ( .A(\ab[10][4] ), .B(n455), .Y(n898) );
  NAND2X1 U1252 ( .A(\SUMB[9][5] ), .B(\ab[10][4] ), .Y(n899) );
  NAND2X1 U1253 ( .A(\SUMB[9][5] ), .B(n455), .Y(n900) );
  NAND3X1 U1254 ( .A(n898), .B(n900), .C(n899), .Y(\CARRYB[10][4] ) );
  NAND2X1 U1255 ( .A(\ab[6][7] ), .B(n679), .Y(n901) );
  NAND2X1 U1256 ( .A(\SUMB[5][8] ), .B(\ab[6][7] ), .Y(n902) );
  NAND2X1 U1257 ( .A(\SUMB[5][8] ), .B(n679), .Y(n903) );
  NAND3X1 U1258 ( .A(n901), .B(n903), .C(n902), .Y(\CARRYB[6][7] ) );
  NAND2X1 U1259 ( .A(\ab[7][6] ), .B(n125), .Y(n904) );
  NAND2X1 U1260 ( .A(\SUMB[6][7] ), .B(\ab[7][6] ), .Y(n905) );
  NAND2X1 U1261 ( .A(\SUMB[6][7] ), .B(n125), .Y(n906) );
  NAND3X1 U1262 ( .A(n904), .B(n905), .C(n906), .Y(\CARRYB[7][6] ) );
  NAND2X1 U1263 ( .A(\ab[9][4] ), .B(n322), .Y(n907) );
  NAND2X1 U1264 ( .A(\SUMB[8][5] ), .B(\ab[9][4] ), .Y(n908) );
  NAND2X1 U1265 ( .A(\SUMB[8][5] ), .B(n322), .Y(n909) );
  NAND3X1 U1266 ( .A(n907), .B(n908), .C(n909), .Y(\CARRYB[9][4] ) );
  NAND2X1 U1267 ( .A(n317), .B(\ab[10][3] ), .Y(n910) );
  NAND2X1 U1268 ( .A(\SUMB[9][4] ), .B(\ab[10][3] ), .Y(n911) );
  NAND2X1 U1269 ( .A(\SUMB[9][4] ), .B(n317), .Y(n912) );
  NAND3X1 U1270 ( .A(n910), .B(n911), .C(n912), .Y(\CARRYB[10][3] ) );
  INVX2 U1271 ( .A(\CARRYB[3][8] ), .Y(n913) );
  NAND2X1 U1272 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .Y(n915) );
  NAND2X1 U1273 ( .A(\SUMB[3][7] ), .B(\ab[4][6] ), .Y(n916) );
  NAND2X1 U1274 ( .A(\SUMB[3][7] ), .B(\CARRYB[3][6] ), .Y(n917) );
  NAND3X1 U1275 ( .A(n915), .B(n916), .C(n917), .Y(\CARRYB[4][6] ) );
  NAND2X1 U1276 ( .A(\ab[5][5] ), .B(n571), .Y(n918) );
  NAND2X1 U1277 ( .A(\SUMB[4][6] ), .B(\ab[5][5] ), .Y(n919) );
  NAND2X1 U1278 ( .A(\SUMB[4][6] ), .B(n571), .Y(n920) );
  NAND3X1 U1279 ( .A(n918), .B(n920), .C(n919), .Y(\CARRYB[5][5] ) );
  NAND2X1 U1280 ( .A(\SUMB[9][3] ), .B(n124), .Y(n921) );
  NAND2X1 U1281 ( .A(\SUMB[9][3] ), .B(\ab[10][2] ), .Y(n922) );
  NAND2X1 U1282 ( .A(n124), .B(\ab[10][2] ), .Y(n923) );
  XOR2X1 U1283 ( .A(n100), .B(n924), .Y(\SUMB[5][6] ) );
  NAND2X1 U1284 ( .A(\ab[4][7] ), .B(n655), .Y(n925) );
  NAND2X1 U1285 ( .A(\SUMB[3][8] ), .B(\ab[4][7] ), .Y(n926) );
  NAND2X1 U1286 ( .A(\SUMB[3][8] ), .B(n655), .Y(n927) );
  NAND3X1 U1287 ( .A(n926), .B(n925), .C(n927), .Y(\CARRYB[4][7] ) );
  NAND2X1 U1288 ( .A(\SUMB[4][7] ), .B(\ab[5][6] ), .Y(n929) );
  NAND2X1 U1289 ( .A(\SUMB[4][7] ), .B(\CARRYB[4][6] ), .Y(n930) );
  NAND3X1 U1290 ( .A(n928), .B(n929), .C(n930), .Y(\CARRYB[5][6] ) );
  NAND2X1 U1291 ( .A(\SUMB[8][4] ), .B(n723), .Y(n931) );
  NAND2X1 U1292 ( .A(\SUMB[8][4] ), .B(\ab[9][3] ), .Y(n932) );
  NAND2X1 U1293 ( .A(n723), .B(\ab[9][3] ), .Y(n933) );
  NAND3X1 U1294 ( .A(n933), .B(n931), .C(n932), .Y(\CARRYB[9][3] ) );
  NAND2X1 U1295 ( .A(n3), .B(\ab[2][8] ), .Y(n934) );
  NAND2X1 U1296 ( .A(\SUMB[1][9] ), .B(\ab[2][8] ), .Y(n935) );
  NAND2X1 U1297 ( .A(\SUMB[1][9] ), .B(n3), .Y(n936) );
  NAND3X1 U1298 ( .A(n934), .B(n935), .C(n936), .Y(\CARRYB[2][8] ) );
  NAND2X1 U1299 ( .A(\ab[3][7] ), .B(n391), .Y(n937) );
  NAND2X1 U1300 ( .A(\SUMB[2][8] ), .B(\ab[3][7] ), .Y(n938) );
  NAND2X1 U1301 ( .A(\SUMB[2][8] ), .B(n391), .Y(n939) );
  NAND3X1 U1302 ( .A(n937), .B(n938), .C(n939), .Y(\CARRYB[3][7] ) );
  NAND2X1 U1303 ( .A(\ab[6][8] ), .B(n946), .Y(n940) );
  NAND2X1 U1304 ( .A(\SUMB[5][9] ), .B(\ab[6][8] ), .Y(n941) );
  NAND2X1 U1305 ( .A(\SUMB[5][9] ), .B(n946), .Y(n942) );
  NAND3X1 U1306 ( .A(n940), .B(n941), .C(n942), .Y(\CARRYB[6][8] ) );
  NAND2X1 U1307 ( .A(n792), .B(\ab[7][7] ), .Y(n943) );
  NAND2X1 U1308 ( .A(\SUMB[6][8] ), .B(\ab[7][7] ), .Y(n944) );
  NAND2X1 U1309 ( .A(\SUMB[6][8] ), .B(n792), .Y(n945) );
  NAND3X1 U1310 ( .A(n944), .B(n943), .C(n945), .Y(\CARRYB[7][7] ) );
  NAND2X1 U1311 ( .A(\ab[2][5] ), .B(n439), .Y(n948) );
  NAND2X1 U1312 ( .A(\ab[2][5] ), .B(\SUMB[1][6] ), .Y(n949) );
  NAND2X1 U1313 ( .A(n439), .B(\SUMB[1][6] ), .Y(n950) );
  NAND3X1 U1314 ( .A(n948), .B(n949), .C(n950), .Y(\CARRYB[2][5] ) );
  NAND2X1 U1315 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .Y(n951) );
  NAND2X1 U1316 ( .A(\ab[3][4] ), .B(\SUMB[2][5] ), .Y(n952) );
  NAND2X1 U1317 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n953) );
  NAND3X1 U1318 ( .A(n951), .B(n952), .C(n953), .Y(\CARRYB[3][4] ) );
  XNOR2X1 U1319 ( .A(\CARRYB[14][0] ), .B(\ab[15][0] ), .Y(n954) );
  XOR2X1 U1320 ( .A(\CARRYB[7][7] ), .B(\ab[8][7] ), .Y(n955) );
  XOR2X1 U1321 ( .A(\SUMB[7][8] ), .B(n955), .Y(\SUMB[8][7] ) );
  NAND2X1 U1322 ( .A(\ab[8][7] ), .B(n969), .Y(n957) );
  NAND2X1 U1323 ( .A(\SUMB[7][8] ), .B(\ab[8][7] ), .Y(n958) );
  NAND2X1 U1324 ( .A(\SUMB[7][8] ), .B(n969), .Y(n959) );
  NAND3X1 U1325 ( .A(n957), .B(n958), .C(n959), .Y(\CARRYB[8][7] ) );
  NAND2X1 U1326 ( .A(\ab[9][6] ), .B(n130), .Y(n960) );
  NAND2X1 U1327 ( .A(\SUMB[8][7] ), .B(\ab[9][6] ), .Y(n961) );
  NAND2X1 U1328 ( .A(n130), .B(\SUMB[8][7] ), .Y(n962) );
  NAND3X1 U1329 ( .A(n960), .B(n961), .C(n962), .Y(\CARRYB[9][6] ) );
  NAND2X1 U1330 ( .A(\ab[14][1] ), .B(n1031), .Y(n963) );
  NAND2X1 U1331 ( .A(\SUMB[13][2] ), .B(\ab[14][1] ), .Y(n964) );
  NAND2X1 U1332 ( .A(\SUMB[13][2] ), .B(n1031), .Y(n965) );
  NAND3X1 U1333 ( .A(n965), .B(n963), .C(n964), .Y(\CARRYB[14][1] ) );
  NAND2X1 U1334 ( .A(n418), .B(\ab[15][0] ), .Y(n966) );
  NAND2X1 U1335 ( .A(\ab[15][0] ), .B(\SUMB[14][1] ), .Y(n967) );
  NAND2X1 U1336 ( .A(n418), .B(\SUMB[14][1] ), .Y(n968) );
  NAND3X1 U1337 ( .A(n966), .B(n968), .C(n967), .Y(\CARRYB[15][0] ) );
  NAND2X1 U1338 ( .A(\CARRYB[6][4] ), .B(\ab[7][4] ), .Y(n970) );
  NAND2X1 U1339 ( .A(\SUMB[6][5] ), .B(\ab[7][4] ), .Y(n971) );
  NAND2X1 U1340 ( .A(\SUMB[6][5] ), .B(n420), .Y(n972) );
  NAND3X1 U1341 ( .A(n970), .B(n971), .C(n972), .Y(\CARRYB[7][4] ) );
  NAND2X1 U1342 ( .A(\ab[8][3] ), .B(n141), .Y(n973) );
  NAND2X1 U1343 ( .A(\SUMB[7][4] ), .B(\ab[8][3] ), .Y(n974) );
  NAND2X1 U1344 ( .A(n348), .B(\SUMB[7][4] ), .Y(n975) );
  NAND3X1 U1345 ( .A(n18), .B(n974), .C(n975), .Y(\CARRYB[8][3] ) );
  XOR2X1 U1346 ( .A(n210), .B(\ab[2][6] ), .Y(n976) );
  NAND2X1 U1347 ( .A(n210), .B(\ab[2][6] ), .Y(n977) );
  NAND2X1 U1348 ( .A(\ab[2][6] ), .B(\SUMB[1][7] ), .Y(n978) );
  NAND2X1 U1349 ( .A(n210), .B(\SUMB[1][7] ), .Y(n979) );
  NAND3X1 U1350 ( .A(n977), .B(n978), .C(n979), .Y(\CARRYB[2][6] ) );
  NAND2X1 U1351 ( .A(\ab[3][5] ), .B(n986), .Y(n980) );
  NAND2X1 U1352 ( .A(\SUMB[2][6] ), .B(\ab[3][5] ), .Y(n981) );
  NAND2X1 U1353 ( .A(\SUMB[2][6] ), .B(n986), .Y(n982) );
  NAND3X1 U1354 ( .A(n980), .B(n981), .C(n982), .Y(\CARRYB[3][5] ) );
  INVX2 U1355 ( .A(\CARRYB[2][5] ), .Y(n985) );
  XOR2X1 U1356 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .Y(n987) );
  XOR2X1 U1357 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .Y(n988) );
  XOR2X1 U1358 ( .A(n988), .B(n476), .Y(\SUMB[4][2] ) );
  NAND2X1 U1359 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .Y(n989) );
  NAND2X1 U1360 ( .A(\ab[3][3] ), .B(\SUMB[2][4] ), .Y(n990) );
  NAND2X1 U1361 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n991) );
  NAND3X1 U1362 ( .A(n989), .B(n990), .C(n991), .Y(\CARRYB[3][3] ) );
  NAND2X1 U1363 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .Y(n992) );
  NAND2X1 U1364 ( .A(\ab[4][2] ), .B(\SUMB[3][3] ), .Y(n993) );
  NAND2X1 U1365 ( .A(\CARRYB[3][2] ), .B(\SUMB[3][3] ), .Y(n994) );
  NAND3X1 U1366 ( .A(n992), .B(n993), .C(n994), .Y(\CARRYB[4][2] ) );
  XOR2X1 U1367 ( .A(n427), .B(\ab[7][1] ), .Y(n995) );
  XOR2X1 U1368 ( .A(n995), .B(n1003), .Y(\SUMB[7][1] ) );
  XOR2X1 U1369 ( .A(\ab[8][0] ), .B(n140), .Y(n996) );
  XOR2X1 U1370 ( .A(n996), .B(\SUMB[7][1] ), .Y(\A1[6] ) );
  NAND2X1 U1371 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .Y(n997) );
  NAND2X1 U1372 ( .A(\ab[7][1] ), .B(\SUMB[6][2] ), .Y(n998) );
  NAND2X1 U1373 ( .A(\SUMB[6][2] ), .B(\CARRYB[6][1] ), .Y(n999) );
  NAND3X1 U1374 ( .A(n998), .B(n997), .C(n999), .Y(\CARRYB[7][1] ) );
  NAND2X1 U1375 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .Y(n1000) );
  NAND2X1 U1376 ( .A(\ab[8][0] ), .B(\SUMB[7][1] ), .Y(n1001) );
  NAND2X1 U1377 ( .A(\CARRYB[7][0] ), .B(\SUMB[7][1] ), .Y(n1002) );
  NAND3X1 U1378 ( .A(n1002), .B(n1001), .C(n1000), .Y(\CARRYB[8][0] ) );
  BUFX2 U1379 ( .A(\SUMB[6][2] ), .Y(n1003) );
  XOR2X1 U1380 ( .A(\CARRYB[2][2] ), .B(\ab[3][2] ), .Y(n1004) );
  XOR2X1 U1381 ( .A(n624), .B(n1004), .Y(\SUMB[3][2] ) );
  NAND2X1 U1382 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(n1005) );
  NAND2X1 U1383 ( .A(\SUMB[2][3] ), .B(\ab[3][2] ), .Y(n1006) );
  NAND2X1 U1384 ( .A(\CARRYB[2][2] ), .B(\ab[3][2] ), .Y(n1007) );
  NAND3X1 U1385 ( .A(n1006), .B(n1005), .C(n1007), .Y(\CARRYB[3][2] ) );
  NAND2X1 U1386 ( .A(\SUMB[6][3] ), .B(\ab[7][2] ), .Y(n1009) );
  NAND2X1 U1387 ( .A(n5), .B(\SUMB[6][3] ), .Y(n1010) );
  NAND3X1 U1388 ( .A(n423), .B(n1009), .C(n1010), .Y(\CARRYB[7][2] ) );
  NAND2X1 U1389 ( .A(\CARRYB[7][1] ), .B(\ab[8][1] ), .Y(n1011) );
  NAND2X1 U1390 ( .A(\SUMB[7][2] ), .B(\ab[8][1] ), .Y(n1012) );
  NAND2X1 U1391 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(n1013) );
  NAND3X1 U1392 ( .A(n1011), .B(n1012), .C(n1013), .Y(\CARRYB[8][1] ) );
  INVX4 U1393 ( .A(A[0]), .Y(n1061) );
  AND2X2 U1394 ( .A(\SUMB[15][1] ), .B(n115), .Y(n1014) );
  AND2X2 U1395 ( .A(\SUMB[15][2] ), .B(\CARRYB[15][1] ), .Y(n1015) );
  AND2X2 U1396 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n1020) );
  INVX1 U1397 ( .A(B[1]), .Y(n1034) );
  INVX2 U1398 ( .A(B[10]), .Y(n1051) );
  INVX2 U1399 ( .A(A[13]), .Y(n1098) );
  INVX2 U1400 ( .A(ZA), .Y(n1096) );
  INVX2 U1401 ( .A(A[14]), .Y(n1097) );
  INVX2 U1402 ( .A(A[4]), .Y(n1068) );
  INVX2 U1403 ( .A(A[5]), .Y(n1070) );
  INVX2 U1404 ( .A(A[6]), .Y(n1072) );
  INVX2 U1405 ( .A(A[7]), .Y(n1074) );
  INVX2 U1406 ( .A(A[9]), .Y(n1078) );
  INVX2 U1407 ( .A(A[8]), .Y(n1076) );
  INVX2 U1408 ( .A(A[10]), .Y(n1080) );
  XOR2X1 U1409 ( .A(\SUMB[15][2] ), .B(\CARRYB[15][1] ), .Y(\A1[15] ) );
  XOR2X1 U1410 ( .A(\SUMB[15][3] ), .B(\CARRYB[15][2] ), .Y(\A1[16] ) );
  XOR2X1 U1411 ( .A(\SUMB[15][4] ), .B(\CARRYB[15][3] ), .Y(\A1[17] ) );
  XOR2X1 U1412 ( .A(\SUMB[15][5] ), .B(\CARRYB[15][4] ), .Y(\A1[18] ) );
  NAND2X1 U1413 ( .A(\SUMB[15][7] ), .B(\CARRYB[15][6] ), .Y(n1023) );
  INVX2 U1414 ( .A(n1023), .Y(\A2[21] ) );
  XOR2X1 U1415 ( .A(\SUMB[15][8] ), .B(\CARRYB[15][7] ), .Y(\A1[21] ) );
  XOR2X1 U1416 ( .A(\SUMB[15][9] ), .B(\CARRYB[15][8] ), .Y(\A1[22] ) );
  XOR2X1 U1417 ( .A(\SUMB[15][10] ), .B(\CARRYB[15][9] ), .Y(\A1[23] ) );
  XOR2X1 U1418 ( .A(\SUMB[15][11] ), .B(\CARRYB[15][10] ), .Y(\A1[24] ) );
  XOR2X1 U1419 ( .A(\SUMB[15][12] ), .B(\CARRYB[15][11] ), .Y(\A1[25] ) );
  XOR2X1 U1420 ( .A(\SUMB[15][13] ), .B(\CARRYB[15][12] ), .Y(\A1[26] ) );
  XOR2X1 U1421 ( .A(\SUMB[15][14] ), .B(\CARRYB[15][13] ), .Y(\A1[27] ) );
  XOR2X1 U1422 ( .A(\SUMB[15][15] ), .B(\CARRYB[15][14] ), .Y(\A1[28] ) );
  XOR2X1 U1423 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U1424 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U1425 ( .A(n1022), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U1426 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U1427 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U1428 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U1429 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(\SUMB[1][10] ) );
  NAND2X1 U1430 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(n1024) );
  XOR2X1 U1431 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(\SUMB[1][11] ) );
  XOR2X1 U1432 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Y(\SUMB[1][12] ) );
  XOR2X1 U1433 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Y(\SUMB[1][13] ) );
  NAND2X1 U1434 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Y(n1025) );
  INVX2 U1435 ( .A(n1025), .Y(\CARRYB[1][13] ) );
  XOR2X1 U1436 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Y(\SUMB[1][14] ) );
  BUFX4 U1437 ( .A(\CARRYB[9][1] ), .Y(n1026) );
  INVX1 U1438 ( .A(n1039), .Y(n1091) );
  INVX1 U1439 ( .A(n1035), .Y(n1093) );
  INVX2 U1440 ( .A(\CARRYB[6][2] ), .Y(n1027) );
  INVX1 U1441 ( .A(n1041), .Y(n1090) );
  INVX4 U1442 ( .A(B[4]), .Y(n1040) );
  INVX2 U1443 ( .A(\CARRYB[10][3] ), .Y(n1028) );
  INVX4 U1444 ( .A(B[2]), .Y(n1036) );
  INVX2 U1445 ( .A(\CARRYB[13][1] ), .Y(n1030) );
  INVX8 U1446 ( .A(n1032), .Y(n1033) );
  INVX8 U1447 ( .A(n1036), .Y(n1037) );
  INVX8 U1448 ( .A(n1038), .Y(n1039) );
  INVX8 U1449 ( .A(n1040), .Y(n1041) );
  INVX8 U1450 ( .A(n1042), .Y(n1043) );
  INVX8 U1451 ( .A(n1044), .Y(n1045) );
  INVX8 U1452 ( .A(n1051), .Y(n1052) );
  INVX8 U1453 ( .A(n1055), .Y(n1056) );
  INVX8 U1454 ( .A(n1057), .Y(n1058) );
  INVX8 U1455 ( .A(n1059), .Y(n1060) );
  INVX8 U1456 ( .A(n1064), .Y(n1065) );
  INVX8 U1457 ( .A(n1066), .Y(n1067) );
  INVX8 U1458 ( .A(n1068), .Y(n1069) );
  INVX8 U1459 ( .A(n1070), .Y(n1071) );
  INVX8 U1460 ( .A(n1072), .Y(n1073) );
  INVX8 U1461 ( .A(n1074), .Y(n1075) );
  INVX8 U1462 ( .A(n1076), .Y(n1077) );
  INVX8 U1463 ( .A(n1078), .Y(n1079) );
  AND2X2 U1464 ( .A(n42), .B(n1060), .Y(\ab[1][14] ) );
  AND2X2 U1465 ( .A(n1060), .B(n103), .Y(\ab[0][14] ) );
  AND2X2 U1466 ( .A(n983), .B(n1058), .Y(\ab[1][13] ) );
  AND2X2 U1467 ( .A(n1058), .B(n1062), .Y(\ab[0][13] ) );
  AND2X2 U1468 ( .A(n42), .B(n1056), .Y(\ab[1][12] ) );
  AND2X2 U1469 ( .A(n1056), .B(n298), .Y(\ab[0][12] ) );
  AND2X2 U1470 ( .A(n42), .B(B[11]), .Y(\ab[1][11] ) );
  AND2X2 U1471 ( .A(n1062), .B(B[11]), .Y(\ab[0][11] ) );
  AND2X2 U1472 ( .A(n983), .B(n1052), .Y(\ab[1][10] ) );
  AND2X2 U1473 ( .A(n1052), .B(n298), .Y(\ab[0][10] ) );
  AND2X2 U1474 ( .A(B[7]), .B(n1062), .Y(\ab[0][7] ) );
  AND2X2 U1475 ( .A(n983), .B(n1043), .Y(\ab[1][5] ) );
  AND2X2 U1476 ( .A(n1043), .B(n103), .Y(\ab[0][5] ) );
  AND2X2 U1477 ( .A(n1041), .B(n983), .Y(\ab[1][4] ) );
  AND2X2 U1478 ( .A(n1041), .B(n103), .Y(\ab[0][4] ) );
  AND2X2 U1479 ( .A(n1039), .B(n984), .Y(\ab[1][3] ) );
  AND2X2 U1480 ( .A(n1039), .B(n105), .Y(\ab[0][3] ) );
  AND2X2 U1481 ( .A(n1037), .B(n894), .Y(\ab[0][2] ) );
  AND2X2 U1482 ( .A(B[1]), .B(n894), .Y(\ab[0][1] ) );
  AND2X2 U1483 ( .A(n984), .B(B[0]), .Y(\ab[1][0] ) );
  AND2X2 U1484 ( .A(n1065), .B(n1060), .Y(\ab[2][14] ) );
  NOR2X1 U1485 ( .A(n984), .B(n1095), .Y(\ab[1][15] ) );
  AND2X2 U1486 ( .A(n1065), .B(n1058), .Y(\ab[2][13] ) );
  AND2X2 U1487 ( .A(n1065), .B(n1056), .Y(\ab[2][12] ) );
  AND2X2 U1488 ( .A(n1065), .B(B[11]), .Y(\ab[2][11] ) );
  AND2X2 U1489 ( .A(n1065), .B(n1052), .Y(\ab[2][10] ) );
  AND2X2 U1490 ( .A(n1065), .B(n579), .Y(\ab[2][9] ) );
  AND2X2 U1491 ( .A(n1065), .B(n529), .Y(\ab[2][8] ) );
  AND2X2 U1492 ( .A(n1065), .B(B[7]), .Y(\ab[2][7] ) );
  AND2X2 U1493 ( .A(n1065), .B(n1045), .Y(\ab[2][6] ) );
  AND2X2 U1494 ( .A(n1065), .B(n1043), .Y(\ab[2][5] ) );
  AND2X2 U1495 ( .A(n1065), .B(n1041), .Y(\ab[2][4] ) );
  AND2X2 U1496 ( .A(n1065), .B(n1039), .Y(\ab[2][3] ) );
  AND2X2 U1497 ( .A(n1065), .B(n1037), .Y(\ab[2][2] ) );
  AND2X2 U1498 ( .A(n153), .B(B[1]), .Y(\ab[2][1] ) );
  AND2X2 U1499 ( .A(n153), .B(n1033), .Y(\ab[2][0] ) );
  AND2X2 U1500 ( .A(n1067), .B(n1060), .Y(\ab[3][14] ) );
  NOR2X1 U1501 ( .A(n153), .B(n1095), .Y(\ab[2][15] ) );
  AND2X2 U1502 ( .A(n1067), .B(n1058), .Y(\ab[3][13] ) );
  AND2X2 U1503 ( .A(n1067), .B(n1056), .Y(\ab[3][12] ) );
  AND2X2 U1504 ( .A(n1067), .B(B[11]), .Y(\ab[3][11] ) );
  AND2X2 U1505 ( .A(n1067), .B(n1052), .Y(\ab[3][10] ) );
  AND2X2 U1506 ( .A(n1067), .B(n579), .Y(\ab[3][9] ) );
  AND2X2 U1507 ( .A(n1067), .B(n529), .Y(\ab[3][8] ) );
  AND2X2 U1508 ( .A(n1067), .B(n1047), .Y(\ab[3][7] ) );
  AND2X2 U1509 ( .A(n1067), .B(n1045), .Y(\ab[3][6] ) );
  AND2X2 U1510 ( .A(n1067), .B(n1043), .Y(\ab[3][5] ) );
  AND2X2 U1511 ( .A(n1067), .B(n1041), .Y(\ab[3][4] ) );
  AND2X2 U1512 ( .A(n1067), .B(n1039), .Y(\ab[3][3] ) );
  AND2X2 U1513 ( .A(n1067), .B(n1037), .Y(\ab[3][2] ) );
  AND2X2 U1514 ( .A(n1067), .B(B[1]), .Y(\ab[3][1] ) );
  AND2X2 U1515 ( .A(n1067), .B(n1033), .Y(\ab[3][0] ) );
  AND2X2 U1516 ( .A(n1069), .B(n1060), .Y(\ab[4][14] ) );
  NOR2X1 U1517 ( .A(n1067), .B(n1095), .Y(\ab[3][15] ) );
  AND2X2 U1518 ( .A(n1069), .B(n1058), .Y(\ab[4][13] ) );
  AND2X2 U1519 ( .A(n1069), .B(n1056), .Y(\ab[4][12] ) );
  AND2X2 U1520 ( .A(n1069), .B(n1054), .Y(\ab[4][11] ) );
  AND2X2 U1521 ( .A(n1069), .B(n1052), .Y(\ab[4][10] ) );
  AND2X2 U1522 ( .A(n1069), .B(n579), .Y(\ab[4][9] ) );
  AND2X2 U1523 ( .A(n1069), .B(n529), .Y(\ab[4][8] ) );
  AND2X2 U1524 ( .A(n1069), .B(n1047), .Y(\ab[4][7] ) );
  AND2X2 U1525 ( .A(n1069), .B(n1045), .Y(\ab[4][6] ) );
  AND2X2 U1526 ( .A(n1069), .B(n1043), .Y(\ab[4][5] ) );
  AND2X2 U1527 ( .A(n1069), .B(n1041), .Y(\ab[4][4] ) );
  AND2X2 U1528 ( .A(n1069), .B(n1039), .Y(\ab[4][3] ) );
  AND2X2 U1529 ( .A(n1069), .B(n1037), .Y(\ab[4][2] ) );
  AND2X2 U1530 ( .A(n1069), .B(n1035), .Y(\ab[4][1] ) );
  AND2X2 U1531 ( .A(n1069), .B(n1033), .Y(\ab[4][0] ) );
  AND2X2 U1532 ( .A(n1071), .B(n1060), .Y(\ab[5][14] ) );
  NOR2X1 U1533 ( .A(n1069), .B(n1095), .Y(\ab[4][15] ) );
  AND2X2 U1534 ( .A(n1071), .B(n1058), .Y(\ab[5][13] ) );
  AND2X2 U1535 ( .A(n1071), .B(n1056), .Y(\ab[5][12] ) );
  AND2X2 U1536 ( .A(n1071), .B(n1054), .Y(\ab[5][11] ) );
  AND2X2 U1537 ( .A(n1071), .B(n1052), .Y(\ab[5][10] ) );
  AND2X2 U1538 ( .A(n1071), .B(n579), .Y(\ab[5][9] ) );
  AND2X2 U1539 ( .A(n1071), .B(n529), .Y(\ab[5][8] ) );
  AND2X2 U1540 ( .A(n1071), .B(n1047), .Y(\ab[5][7] ) );
  AND2X2 U1541 ( .A(n1071), .B(n1045), .Y(\ab[5][6] ) );
  AND2X2 U1542 ( .A(n1071), .B(n1043), .Y(\ab[5][5] ) );
  AND2X2 U1543 ( .A(n1071), .B(n1041), .Y(\ab[5][4] ) );
  AND2X2 U1544 ( .A(n1071), .B(n1039), .Y(\ab[5][3] ) );
  AND2X2 U1545 ( .A(n1071), .B(n1037), .Y(\ab[5][2] ) );
  AND2X2 U1546 ( .A(n1071), .B(n1035), .Y(\ab[5][1] ) );
  AND2X2 U1547 ( .A(n1071), .B(n1033), .Y(\ab[5][0] ) );
  AND2X2 U1548 ( .A(n1073), .B(n1060), .Y(\ab[6][14] ) );
  NOR2X1 U1549 ( .A(n1071), .B(n1095), .Y(\ab[5][15] ) );
  AND2X2 U1550 ( .A(n1073), .B(n1058), .Y(\ab[6][13] ) );
  AND2X2 U1551 ( .A(n1073), .B(n1056), .Y(\ab[6][12] ) );
  AND2X2 U1552 ( .A(n1073), .B(n1054), .Y(\ab[6][11] ) );
  AND2X2 U1553 ( .A(n1073), .B(n1052), .Y(\ab[6][10] ) );
  AND2X2 U1554 ( .A(n1073), .B(n579), .Y(\ab[6][9] ) );
  AND2X2 U1555 ( .A(n1073), .B(n529), .Y(\ab[6][8] ) );
  AND2X2 U1556 ( .A(n1073), .B(n1047), .Y(\ab[6][7] ) );
  AND2X2 U1557 ( .A(n1073), .B(n1045), .Y(\ab[6][6] ) );
  AND2X2 U1558 ( .A(n1073), .B(n1043), .Y(\ab[6][5] ) );
  AND2X2 U1559 ( .A(n1073), .B(n1041), .Y(\ab[6][4] ) );
  AND2X2 U1560 ( .A(n1073), .B(n1039), .Y(\ab[6][3] ) );
  AND2X2 U1561 ( .A(n1073), .B(n1037), .Y(\ab[6][2] ) );
  AND2X2 U1562 ( .A(n1073), .B(n1035), .Y(\ab[6][1] ) );
  AND2X2 U1563 ( .A(n1073), .B(n1033), .Y(\ab[6][0] ) );
  AND2X2 U1564 ( .A(n1075), .B(n1060), .Y(\ab[7][14] ) );
  NOR2X1 U1565 ( .A(n1073), .B(n1095), .Y(\ab[6][15] ) );
  AND2X2 U1566 ( .A(n1075), .B(n1058), .Y(\ab[7][13] ) );
  AND2X2 U1567 ( .A(n1075), .B(n1056), .Y(\ab[7][12] ) );
  AND2X2 U1568 ( .A(n1075), .B(n1054), .Y(\ab[7][11] ) );
  AND2X2 U1569 ( .A(n1075), .B(n1052), .Y(\ab[7][10] ) );
  AND2X2 U1570 ( .A(n1075), .B(n579), .Y(\ab[7][9] ) );
  AND2X2 U1571 ( .A(n1075), .B(n529), .Y(\ab[7][8] ) );
  AND2X2 U1572 ( .A(n1075), .B(n1047), .Y(\ab[7][7] ) );
  AND2X2 U1573 ( .A(n1075), .B(n1045), .Y(\ab[7][6] ) );
  AND2X2 U1574 ( .A(n1075), .B(n1043), .Y(\ab[7][5] ) );
  AND2X2 U1575 ( .A(n1075), .B(n1041), .Y(\ab[7][4] ) );
  AND2X2 U1576 ( .A(n1075), .B(n1039), .Y(\ab[7][3] ) );
  AND2X2 U1577 ( .A(n1075), .B(n1037), .Y(\ab[7][2] ) );
  AND2X2 U1578 ( .A(n1075), .B(n1035), .Y(\ab[7][1] ) );
  AND2X2 U1579 ( .A(n1075), .B(n1033), .Y(\ab[7][0] ) );
  AND2X2 U1580 ( .A(n1077), .B(n1060), .Y(\ab[8][14] ) );
  NOR2X1 U1581 ( .A(n1075), .B(n1095), .Y(\ab[7][15] ) );
  AND2X2 U1582 ( .A(n1077), .B(n1058), .Y(\ab[8][13] ) );
  AND2X2 U1583 ( .A(n1077), .B(n1056), .Y(\ab[8][12] ) );
  AND2X2 U1584 ( .A(n1077), .B(n1054), .Y(\ab[8][11] ) );
  AND2X2 U1585 ( .A(n1077), .B(n1052), .Y(\ab[8][10] ) );
  AND2X2 U1586 ( .A(n1077), .B(n579), .Y(\ab[8][9] ) );
  AND2X2 U1587 ( .A(n1077), .B(n529), .Y(\ab[8][8] ) );
  AND2X2 U1588 ( .A(n1077), .B(n1047), .Y(\ab[8][7] ) );
  AND2X2 U1589 ( .A(n1077), .B(n1045), .Y(\ab[8][6] ) );
  AND2X2 U1590 ( .A(n1077), .B(n1043), .Y(\ab[8][5] ) );
  AND2X2 U1591 ( .A(n1077), .B(n1041), .Y(\ab[8][4] ) );
  AND2X2 U1592 ( .A(n1077), .B(n1039), .Y(\ab[8][3] ) );
  AND2X2 U1593 ( .A(n1077), .B(n1037), .Y(\ab[8][2] ) );
  AND2X2 U1594 ( .A(n1077), .B(n1035), .Y(\ab[8][1] ) );
  AND2X2 U1595 ( .A(n1077), .B(n1033), .Y(\ab[8][0] ) );
  AND2X2 U1596 ( .A(n1079), .B(n1060), .Y(\ab[9][14] ) );
  NOR2X1 U1597 ( .A(n1077), .B(n1095), .Y(\ab[8][15] ) );
  AND2X2 U1598 ( .A(n1079), .B(n1058), .Y(\ab[9][13] ) );
  AND2X2 U1599 ( .A(n1079), .B(n1056), .Y(\ab[9][12] ) );
  AND2X2 U1600 ( .A(n1079), .B(n1054), .Y(\ab[9][11] ) );
  AND2X2 U1601 ( .A(n1079), .B(n1052), .Y(\ab[9][10] ) );
  AND2X2 U1602 ( .A(n1079), .B(n579), .Y(\ab[9][9] ) );
  AND2X2 U1603 ( .A(n1079), .B(n529), .Y(\ab[9][8] ) );
  AND2X2 U1604 ( .A(n1079), .B(n1047), .Y(\ab[9][7] ) );
  AND2X2 U1605 ( .A(n1079), .B(n1045), .Y(\ab[9][6] ) );
  AND2X2 U1606 ( .A(n1079), .B(n1043), .Y(\ab[9][5] ) );
  AND2X2 U1607 ( .A(n1079), .B(n1041), .Y(\ab[9][4] ) );
  AND2X2 U1608 ( .A(n1079), .B(n1039), .Y(\ab[9][3] ) );
  AND2X2 U1609 ( .A(n1079), .B(n1037), .Y(\ab[9][2] ) );
  AND2X2 U1610 ( .A(n1079), .B(n1035), .Y(\ab[9][1] ) );
  AND2X2 U1611 ( .A(n1079), .B(n1033), .Y(\ab[9][0] ) );
  AND2X2 U1612 ( .A(n1081), .B(n1060), .Y(\ab[10][14] ) );
  NOR2X1 U1613 ( .A(n1079), .B(n1095), .Y(\ab[9][15] ) );
  AND2X2 U1614 ( .A(n1081), .B(n1058), .Y(\ab[10][13] ) );
  AND2X2 U1615 ( .A(n1081), .B(n1056), .Y(\ab[10][12] ) );
  AND2X2 U1616 ( .A(n1081), .B(n1054), .Y(\ab[10][11] ) );
  AND2X2 U1617 ( .A(n1081), .B(n1052), .Y(\ab[10][10] ) );
  AND2X2 U1618 ( .A(n1081), .B(n579), .Y(\ab[10][9] ) );
  AND2X2 U1619 ( .A(n1081), .B(n529), .Y(\ab[10][8] ) );
  AND2X2 U1620 ( .A(n1081), .B(n1047), .Y(\ab[10][7] ) );
  AND2X2 U1621 ( .A(n1081), .B(n1045), .Y(\ab[10][6] ) );
  AND2X2 U1622 ( .A(n1081), .B(n1043), .Y(\ab[10][5] ) );
  AND2X2 U1623 ( .A(n1081), .B(n1041), .Y(\ab[10][4] ) );
  AND2X2 U1624 ( .A(n1081), .B(n1039), .Y(\ab[10][3] ) );
  AND2X2 U1625 ( .A(n1081), .B(n1037), .Y(\ab[10][2] ) );
  AND2X2 U1626 ( .A(n1081), .B(n1035), .Y(\ab[10][1] ) );
  AND2X2 U1627 ( .A(n1081), .B(n1033), .Y(\ab[10][0] ) );
  AND2X2 U1628 ( .A(A[11]), .B(n1060), .Y(\ab[11][14] ) );
  NOR2X1 U1629 ( .A(n1081), .B(n1095), .Y(\ab[10][15] ) );
  AND2X2 U1630 ( .A(A[11]), .B(n1058), .Y(\ab[11][13] ) );
  AND2X2 U1631 ( .A(A[11]), .B(n1056), .Y(\ab[11][12] ) );
  AND2X2 U1632 ( .A(A[11]), .B(n1054), .Y(\ab[11][11] ) );
  AND2X2 U1633 ( .A(A[11]), .B(n1052), .Y(\ab[11][10] ) );
  AND2X2 U1634 ( .A(A[11]), .B(n579), .Y(\ab[11][9] ) );
  AND2X2 U1635 ( .A(A[11]), .B(n529), .Y(\ab[11][8] ) );
  AND2X2 U1636 ( .A(A[11]), .B(n1047), .Y(\ab[11][7] ) );
  AND2X2 U1637 ( .A(A[11]), .B(n1045), .Y(\ab[11][6] ) );
  AND2X2 U1638 ( .A(A[11]), .B(n1043), .Y(\ab[11][5] ) );
  AND2X2 U1639 ( .A(A[11]), .B(n1041), .Y(\ab[11][4] ) );
  AND2X2 U1640 ( .A(A[11]), .B(n1039), .Y(\ab[11][3] ) );
  AND2X2 U1641 ( .A(A[11]), .B(n1037), .Y(\ab[11][2] ) );
  AND2X2 U1642 ( .A(A[11]), .B(n1035), .Y(\ab[11][1] ) );
  AND2X2 U1643 ( .A(A[11]), .B(n1033), .Y(\ab[11][0] ) );
  AND2X2 U1644 ( .A(A[12]), .B(n1060), .Y(\ab[12][14] ) );
  NOR2X1 U1645 ( .A(A[11]), .B(n1095), .Y(\ab[11][15] ) );
  AND2X2 U1646 ( .A(A[12]), .B(n1058), .Y(\ab[12][13] ) );
  AND2X2 U1647 ( .A(A[12]), .B(n1056), .Y(\ab[12][12] ) );
  AND2X2 U1648 ( .A(A[12]), .B(n1054), .Y(\ab[12][11] ) );
  AND2X2 U1649 ( .A(A[12]), .B(n1052), .Y(\ab[12][10] ) );
  AND2X2 U1650 ( .A(A[12]), .B(n579), .Y(\ab[12][9] ) );
  AND2X2 U1651 ( .A(A[12]), .B(n529), .Y(\ab[12][8] ) );
  AND2X2 U1652 ( .A(A[12]), .B(n1047), .Y(\ab[12][7] ) );
  AND2X2 U1653 ( .A(A[12]), .B(n1045), .Y(\ab[12][6] ) );
  AND2X2 U1654 ( .A(A[12]), .B(n1043), .Y(\ab[12][5] ) );
  AND2X2 U1655 ( .A(A[12]), .B(n1041), .Y(\ab[12][4] ) );
  AND2X2 U1656 ( .A(A[12]), .B(n1039), .Y(\ab[12][3] ) );
  AND2X2 U1657 ( .A(A[12]), .B(n1037), .Y(\ab[12][2] ) );
  AND2X2 U1658 ( .A(A[12]), .B(n1035), .Y(\ab[12][1] ) );
  AND2X2 U1659 ( .A(A[12]), .B(n1033), .Y(\ab[12][0] ) );
  NOR2X1 U1660 ( .A(n1098), .B(n1082), .Y(\ab[13][14] ) );
  NOR2X1 U1661 ( .A(A[12]), .B(n1095), .Y(\ab[12][15] ) );
  INVX2 U1662 ( .A(n1058), .Y(n1083) );
  NOR2X1 U1663 ( .A(n1098), .B(n1083), .Y(\ab[13][13] ) );
  NOR2X1 U1664 ( .A(n1098), .B(n1084), .Y(\ab[13][12] ) );
  NOR2X1 U1665 ( .A(n1098), .B(n1053), .Y(\ab[13][11] ) );
  NOR2X1 U1666 ( .A(n1098), .B(n1085), .Y(\ab[13][10] ) );
  NOR2X1 U1667 ( .A(n1098), .B(n1086), .Y(\ab[13][9] ) );
  NOR2X1 U1668 ( .A(n1098), .B(n1048), .Y(\ab[13][8] ) );
  NOR2X1 U1669 ( .A(n1098), .B(n1087), .Y(\ab[13][7] ) );
  NOR2X1 U1670 ( .A(n1098), .B(n1088), .Y(\ab[13][6] ) );
  NOR2X1 U1671 ( .A(n1098), .B(n1089), .Y(\ab[13][5] ) );
  NOR2X1 U1672 ( .A(n1098), .B(n1090), .Y(\ab[13][4] ) );
  NOR2X1 U1673 ( .A(n1098), .B(n1091), .Y(\ab[13][3] ) );
  NOR2X1 U1674 ( .A(n1098), .B(n1092), .Y(\ab[13][2] ) );
  NOR2X1 U1675 ( .A(n1098), .B(n1093), .Y(\ab[13][1] ) );
  NOR2X1 U1676 ( .A(n1098), .B(n1032), .Y(\ab[13][0] ) );
  NOR2X1 U1677 ( .A(n1097), .B(n1082), .Y(\ab[14][14] ) );
  NOR2X1 U1678 ( .A(A[13]), .B(n1095), .Y(\ab[13][15] ) );
  NOR2X1 U1679 ( .A(n1097), .B(n1083), .Y(\ab[14][13] ) );
  NOR2X1 U1680 ( .A(n1097), .B(n1084), .Y(\ab[14][12] ) );
  NOR2X1 U1681 ( .A(n1097), .B(n1053), .Y(\ab[14][11] ) );
  NOR2X1 U1682 ( .A(n1097), .B(n1085), .Y(\ab[14][10] ) );
  NOR2X1 U1683 ( .A(n1097), .B(n1086), .Y(\ab[14][9] ) );
  NOR2X1 U1684 ( .A(n1097), .B(n1048), .Y(\ab[14][8] ) );
  NOR2X1 U1685 ( .A(n1097), .B(n1087), .Y(\ab[14][7] ) );
  NOR2X1 U1686 ( .A(n1097), .B(n1088), .Y(\ab[14][6] ) );
  NOR2X1 U1687 ( .A(n1097), .B(n1089), .Y(\ab[14][5] ) );
  NOR2X1 U1688 ( .A(n1097), .B(n1090), .Y(\ab[14][4] ) );
  NOR2X1 U1689 ( .A(n1097), .B(n1091), .Y(\ab[14][3] ) );
  NOR2X1 U1690 ( .A(n1097), .B(n1092), .Y(\ab[14][2] ) );
  NOR2X1 U1691 ( .A(n1097), .B(n1093), .Y(\ab[14][1] ) );
  NOR2X1 U1692 ( .A(n1097), .B(n1032), .Y(\ab[14][0] ) );
  NOR2X1 U1693 ( .A(n1096), .B(n1095), .Y(\ab[15][15] ) );
  NOR2X1 U1694 ( .A(A[14]), .B(n1095), .Y(\ab[14][15] ) );
  AND2X2 U1695 ( .A(n1033), .B(n894), .Y(PRODUCT[0]) );
  INVX2 U1696 ( .A(\CARRYB[15][15] ), .Y(n1094) );
  NOR2X1 U1697 ( .A(n579), .B(n1096), .Y(\ab[15][9] ) );
  NOR2X1 U1698 ( .A(n529), .B(n1096), .Y(\ab[15][8] ) );
  NOR2X1 U1699 ( .A(n1047), .B(n1096), .Y(\ab[15][7] ) );
  NOR2X1 U1700 ( .A(n1045), .B(n1096), .Y(\ab[15][6] ) );
  NOR2X1 U1701 ( .A(n1043), .B(n1096), .Y(\ab[15][5] ) );
  NOR2X1 U1702 ( .A(n1041), .B(n1096), .Y(\ab[15][4] ) );
  NOR2X1 U1703 ( .A(n1039), .B(n1096), .Y(\ab[15][3] ) );
  NOR2X1 U1704 ( .A(n1037), .B(n1096), .Y(\ab[15][2] ) );
  NOR2X1 U1705 ( .A(n1035), .B(n1096), .Y(\ab[15][1] ) );
  NOR2X1 U1706 ( .A(n1060), .B(n1096), .Y(\ab[15][14] ) );
  NOR2X1 U1707 ( .A(n1058), .B(n1096), .Y(\ab[15][13] ) );
  NOR2X1 U1708 ( .A(n1056), .B(n1096), .Y(\ab[15][12] ) );
  NOR2X1 U1709 ( .A(n1054), .B(n1096), .Y(\ab[15][11] ) );
  NOR2X1 U1710 ( .A(n1052), .B(n1096), .Y(\ab[15][10] ) );
  NOR2X1 U1711 ( .A(n1033), .B(n1096), .Y(\ab[15][0] ) );
endmodule


module matrix_math_DW01_add_24 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] ,
         \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48;
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  OR2X2 U2 ( .A(A[17]), .B(B[17]), .Y(n1) );
  BUFX2 U3 ( .A(A[14]), .Y(n2) );
  BUFX2 U4 ( .A(B[14]), .Y(n3) );
  OR2X1 U5 ( .A(n2), .B(n3), .Y(n43) );
  XOR2X1 U6 ( .A(n4), .B(n24), .Y(SUM[19]) );
  INVX1 U7 ( .A(n22), .Y(n4) );
  OR2X2 U8 ( .A(A[15]), .B(B[15]), .Y(n8) );
  XNOR2X1 U9 ( .A(n38), .B(n5), .Y(SUM[17]) );
  NAND2X1 U10 ( .A(n1), .B(n36), .Y(n5) );
  NOR2X1 U11 ( .A(A[17]), .B(B[17]), .Y(n6) );
  AND2X2 U12 ( .A(n10), .B(n1), .Y(n7) );
  INVX1 U13 ( .A(n39), .Y(n10) );
  OR2X1 U14 ( .A(A[15]), .B(B[15]), .Y(n42) );
  XNOR2X1 U15 ( .A(n9), .B(n44), .Y(SUM[16]) );
  NAND2X1 U16 ( .A(n45), .B(n41), .Y(n9) );
  INVX1 U17 ( .A(n37), .Y(n39) );
  AND2X2 U18 ( .A(A[14]), .B(B[14]), .Y(n46) );
  XOR2X1 U19 ( .A(n14), .B(n11), .Y(SUM[21]) );
  XNOR2X1 U20 ( .A(B[21]), .B(A[21]), .Y(n11) );
  XNOR2X1 U21 ( .A(n32), .B(n33), .Y(SUM[18]) );
  XOR2X1 U22 ( .A(n48), .B(n47), .Y(SUM[15]) );
  AND2X2 U23 ( .A(n40), .B(n41), .Y(n12) );
  AND2X2 U24 ( .A(n43), .B(n48), .Y(SUM[14]) );
  AOI21X1 U25 ( .A(n20), .B(n15), .C(n16), .Y(n14) );
  INVX2 U26 ( .A(n17), .Y(n16) );
  XNOR2X1 U27 ( .A(n21), .B(n20), .Y(SUM[20]) );
  NAND2X1 U28 ( .A(n15), .B(n17), .Y(n21) );
  NAND2X1 U29 ( .A(B[20]), .B(A[20]), .Y(n17) );
  OR2X2 U30 ( .A(A[20]), .B(B[20]), .Y(n15) );
  NAND2X1 U31 ( .A(n19), .B(n18), .Y(n20) );
  NAND2X1 U32 ( .A(n22), .B(n23), .Y(n19) );
  NAND2X1 U33 ( .A(n23), .B(n18), .Y(n24) );
  NAND2X1 U34 ( .A(A[19]), .B(B[19]), .Y(n18) );
  OR2X2 U35 ( .A(A[19]), .B(B[19]), .Y(n23) );
  OAI21X1 U36 ( .A(n12), .B(n25), .C(n26), .Y(n22) );
  AOI21X1 U37 ( .A(n28), .B(n27), .C(n29), .Y(n26) );
  INVX2 U38 ( .A(n30), .Y(n29) );
  NAND2X1 U39 ( .A(n28), .B(n7), .Y(n25) );
  NAND2X1 U40 ( .A(n30), .B(n28), .Y(n33) );
  OR2X2 U41 ( .A(A[18]), .B(B[18]), .Y(n28) );
  NAND2X1 U42 ( .A(B[18]), .B(A[18]), .Y(n30) );
  OAI21X1 U43 ( .A(n12), .B(n31), .C(n34), .Y(n32) );
  INVX2 U44 ( .A(n27), .Y(n34) );
  OAI21X1 U45 ( .A(n6), .B(n35), .C(n36), .Y(n27) );
  NAND2X1 U46 ( .A(n10), .B(n1), .Y(n31) );
  NAND2X1 U47 ( .A(A[17]), .B(B[17]), .Y(n36) );
  OAI21X1 U48 ( .A(n39), .B(n12), .C(n35), .Y(n38) );
  NAND2X1 U49 ( .A(n8), .B(n46), .Y(n40) );
  NAND2X1 U50 ( .A(n35), .B(n37), .Y(n44) );
  NAND2X1 U51 ( .A(A[16]), .B(B[16]), .Y(n35) );
  OR2X2 U52 ( .A(A[16]), .B(B[16]), .Y(n37) );
  NAND2X1 U53 ( .A(n42), .B(n46), .Y(n45) );
  NAND2X1 U54 ( .A(n41), .B(n8), .Y(n47) );
  NAND2X1 U55 ( .A(A[15]), .B(B[15]), .Y(n41) );
  NAND2X1 U56 ( .A(n3), .B(n2), .Y(n48) );
endmodule


module matrix_math_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] ,
         \ab[2][6] , \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] ,
         \ab[2][0] , \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] ,
         \ab[1][11] , \ab[1][10] , \ab[1][8] , \ab[1][6] , \ab[1][5] ,
         \ab[1][3] , \ab[1][1] , \ab[1][0] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][11] , \ab[0][10] , \ab[0][9] , \ab[0][8] ,
         \ab[0][7] , \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] ,
         \ab[0][1] , \CARRYB[15][15] , \CARRYB[15][14] , \CARRYB[15][13] ,
         \CARRYB[15][12] , \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] ,
         \CARRYB[15][8] , \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] ,
         \CARRYB[15][4] , \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] ,
         \CARRYB[15][0] , \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] ,
         \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][14] ,
         \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] ,
         \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] ,
         \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][13] , \CARRYB[1][12] ,
         \CARRYB[1][9] , \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] ,
         \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] ,
         \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] ,
         \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[15][0] , \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] ,
         \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] ,
         \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] ,
         \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][14] ,
         \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] ,
         \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] ,
         \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] ,
         \SUMB[13][1] , \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] ,
         \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] ,
         \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] ,
         \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][14] ,
         \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] ,
         \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][6] , \SUMB[11][5] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] , \SUMB[10][13] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] ,
         \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][10] , \SUMB[2][9] ,
         \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , ZA, ZB,
         \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[14] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;
  assign ZA = A[15];
  assign ZB = B[15];

  FAX1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .C(\SUMB[14][6] ), .YC(
        \CARRYB[15][5] ), .YS(\SUMB[15][5] ) );
  FAX1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .C(\SUMB[14][9] ), .YC(
        \CARRYB[15][8] ), .YS(\SUMB[15][8] ) );
  FAX1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .C(\SUMB[14][10] ), .YC(
        \CARRYB[15][9] ), .YS(\SUMB[15][9] ) );
  FAX1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .C(\SUMB[14][11] ), 
        .YC(\CARRYB[15][10] ), .YS(\SUMB[15][10] ) );
  FAX1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .C(\SUMB[14][12] ), 
        .YC(\CARRYB[15][11] ), .YS(\SUMB[15][11] ) );
  FAX1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .C(\SUMB[14][13] ), 
        .YC(\CARRYB[15][12] ), .YS(\SUMB[15][12] ) );
  FAX1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .C(\SUMB[14][14] ), 
        .YC(\CARRYB[15][13] ), .YS(\SUMB[15][13] ) );
  FAX1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .C(\ab[14][15] ), .YC(
        \CARRYB[15][14] ), .YS(\SUMB[15][14] ) );
  FAX1 S14_15 ( .A(n1050), .B(n1049), .C(\ab[15][15] ), .YC(\CARRYB[15][15] ), 
        .YS(\SUMB[15][15] ) );
  FAX1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .C(\SUMB[13][10] ), 
        .YC(\CARRYB[14][9] ), .YS(\SUMB[14][9] ) );
  FAX1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .C(\SUMB[13][11] ), 
        .YC(\CARRYB[14][10] ), .YS(\SUMB[14][10] ) );
  FAX1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .C(\SUMB[13][12] ), 
        .YC(\CARRYB[14][11] ), .YS(\SUMB[14][11] ) );
  FAX1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .C(\SUMB[13][13] ), 
        .YC(\CARRYB[14][12] ), .YS(\SUMB[14][12] ) );
  FAX1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .C(\SUMB[13][14] ), 
        .YC(\CARRYB[14][13] ), .YS(\SUMB[14][13] ) );
  FAX1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .C(\ab[13][15] ), 
        .YC(\CARRYB[14][14] ), .YS(\SUMB[14][14] ) );
  FAX1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .C(\SUMB[12][10] ), 
        .YC(\CARRYB[13][9] ), .YS(\SUMB[13][9] ) );
  FAX1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .C(\SUMB[12][11] ), 
        .YC(\CARRYB[13][10] ), .YS(\SUMB[13][10] ) );
  FAX1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .C(\SUMB[12][12] ), 
        .YC(\CARRYB[13][11] ), .YS(\SUMB[13][11] ) );
  FAX1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .C(\SUMB[12][13] ), 
        .YC(\CARRYB[13][12] ), .YS(\SUMB[13][12] ) );
  FAX1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .C(\SUMB[12][14] ), 
        .YC(\CARRYB[13][13] ), .YS(\SUMB[13][13] ) );
  FAX1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .C(\ab[12][15] ), 
        .YC(\CARRYB[13][14] ), .YS(\SUMB[13][14] ) );
  FAX1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .C(\SUMB[11][12] ), 
        .YC(\CARRYB[12][11] ), .YS(\SUMB[12][11] ) );
  FAX1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .C(\SUMB[11][13] ), 
        .YC(\CARRYB[12][12] ), .YS(\SUMB[12][12] ) );
  FAX1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .C(\SUMB[11][14] ), 
        .YC(\CARRYB[12][13] ), .YS(\SUMB[12][13] ) );
  FAX1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .C(\ab[11][15] ), 
        .YC(\CARRYB[12][14] ), .YS(\SUMB[12][14] ) );
  FAX1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .C(\SUMB[10][10] ), 
        .YC(\CARRYB[11][9] ), .YS(\SUMB[11][9] ) );
  FAX1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .C(\SUMB[10][12] ), 
        .YC(\CARRYB[11][11] ), .YS(\SUMB[11][11] ) );
  FAX1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .C(\SUMB[10][13] ), 
        .YC(\CARRYB[11][12] ), .YS(\SUMB[11][12] ) );
  FAX1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .C(\SUMB[10][14] ), 
        .YC(\CARRYB[11][13] ), .YS(\SUMB[11][13] ) );
  FAX1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .C(\ab[10][15] ), 
        .YC(\CARRYB[11][14] ), .YS(\SUMB[11][14] ) );
  FAX1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .C(\SUMB[9][11] ), 
        .YC(\CARRYB[10][10] ), .YS(\SUMB[10][10] ) );
  FAX1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .C(\SUMB[9][12] ), 
        .YC(\CARRYB[10][11] ), .YS(\SUMB[10][11] ) );
  FAX1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .C(\SUMB[9][13] ), 
        .YC(\CARRYB[10][12] ), .YS(\SUMB[10][12] ) );
  FAX1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .C(\SUMB[9][14] ), 
        .YC(\CARRYB[10][13] ), .YS(\SUMB[10][13] ) );
  FAX1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .C(\ab[9][15] ), .YC(
        \CARRYB[10][14] ), .YS(\SUMB[10][14] ) );
  FAX1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .C(\SUMB[8][13] ), .YC(
        \CARRYB[9][12] ), .YS(\SUMB[9][12] ) );
  FAX1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .C(\ab[8][15] ), .YC(
        \CARRYB[9][14] ), .YS(\SUMB[9][14] ) );
  FAX1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .C(\SUMB[7][1] ), .YC(
        \CARRYB[8][0] ), .YS(\A1[6] ) );
  FAX1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .C(\SUMB[7][10] ), .YC(
        \CARRYB[8][9] ), .YS(\SUMB[8][9] ) );
  FAX1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .C(\ab[7][15] ), .YC(
        \CARRYB[8][14] ), .YS(\SUMB[8][14] ) );
  FAX1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .C(\SUMB[6][14] ), .YC(
        \CARRYB[7][13] ), .YS(\SUMB[7][13] ) );
  FAX1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .C(\ab[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S1_6_0 ( .A(\ab[6][0] ), .B(\SUMB[5][1] ), .C(\CARRYB[5][0] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S3_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .C(\ab[5][15] ), .YC(
        \CARRYB[6][14] ), .YS(\SUMB[6][14] ) );
  FAX1 S1_5_0 ( .A(\ab[5][0] ), .B(n908), .C(\SUMB[4][1] ), .YC(\CARRYB[5][0] ), .YS(\A1[3] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(n906), .C(\SUMB[3][1] ), .YC(\CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S3_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .C(\ab[3][15] ), .YC(
        \CARRYB[4][14] ), .YS(\SUMB[4][14] ) );
  FAX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(\A1[1] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n74), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n969), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), .YS(\SUMB[2][1] ) );
  matrix_math_DW01_add_24 FS_1 ( .A({n1048, \A1[28] , \A1[27] , \A1[26] , 
        \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , 
        \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n73, n72, n71, n70, 
        n69, n68, n67, n66, n80, n973, n968, n967, n966, n971, n972, \A2[14] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, PRODUCT[23:2]}) );
  XOR2X1 U2 ( .A(n14), .B(n3), .Y(\SUMB[9][5] ) );
  XNOR2X1 U3 ( .A(n129), .B(n130), .Y(n3) );
  XOR2X1 U4 ( .A(n4), .B(n146), .Y(\SUMB[10][5] ) );
  XNOR2X1 U5 ( .A(\CARRYB[9][5] ), .B(n157), .Y(n4) );
  BUFX2 U6 ( .A(n76), .Y(n5) );
  XNOR2X1 U7 ( .A(n6), .B(\SUMB[4][10] ), .Y(\SUMB[5][9] ) );
  XNOR2X1 U8 ( .A(\CARRYB[4][9] ), .B(\ab[5][9] ), .Y(n6) );
  XNOR2X1 U9 ( .A(n7), .B(\SUMB[5][9] ), .Y(\SUMB[6][8] ) );
  XOR2X1 U10 ( .A(\CARRYB[5][8] ), .B(n175), .Y(n7) );
  XNOR2X1 U11 ( .A(n8), .B(n297), .Y(n223) );
  XOR2X1 U12 ( .A(n222), .B(n82), .Y(n8) );
  INVX2 U13 ( .A(n763), .Y(n9) );
  INVX2 U14 ( .A(n9), .Y(n10) );
  BUFX2 U15 ( .A(n606), .Y(n11) );
  BUFX2 U16 ( .A(n639), .Y(n12) );
  INVX2 U17 ( .A(\SUMB[9][9] ), .Y(n59) );
  BUFX2 U18 ( .A(n765), .Y(n13) );
  XOR2X1 U19 ( .A(\CARRYB[8][5] ), .B(n224), .Y(n14) );
  BUFX2 U20 ( .A(\CARRYB[5][3] ), .Y(n15) );
  NAND3X1 U21 ( .A(n735), .B(n734), .C(n733), .Y(n16) );
  INVX2 U22 ( .A(\SUMB[12][2] ), .Y(n320) );
  XNOR2X1 U23 ( .A(n17), .B(\SUMB[14][1] ), .Y(\SUMB[15][0] ) );
  XNOR2X1 U24 ( .A(\CARRYB[14][0] ), .B(n50), .Y(n17) );
  XNOR2X1 U25 ( .A(n18), .B(n253), .Y(\SUMB[9][4] ) );
  XOR2X1 U26 ( .A(\CARRYB[8][4] ), .B(\ab[9][4] ), .Y(n18) );
  BUFX2 U27 ( .A(\CARRYB[12][7] ), .Y(n19) );
  XOR2X1 U28 ( .A(\SUMB[8][7] ), .B(n20), .Y(\SUMB[9][6] ) );
  XOR2X1 U29 ( .A(\CARRYB[8][6] ), .B(\ab[9][6] ), .Y(n20) );
  BUFX2 U30 ( .A(\SUMB[15][3] ), .Y(n21) );
  AND2X2 U31 ( .A(\CARRYB[15][2] ), .B(n21), .Y(n966) );
  XOR2X1 U32 ( .A(n22), .B(\SUMB[8][8] ), .Y(\SUMB[9][7] ) );
  XOR2X1 U33 ( .A(\CARRYB[8][7] ), .B(\ab[9][7] ), .Y(n22) );
  XOR2X1 U34 ( .A(n23), .B(n5), .Y(\SUMB[12][6] ) );
  XNOR2X1 U35 ( .A(\CARRYB[11][6] ), .B(n244), .Y(n23) );
  BUFX2 U36 ( .A(n898), .Y(n24) );
  XOR2X1 U37 ( .A(\CARRYB[11][4] ), .B(n25), .Y(n339) );
  INVX8 U38 ( .A(\ab[12][4] ), .Y(n25) );
  BUFX2 U39 ( .A(\CARRYB[7][11] ), .Y(n26) );
  INVX2 U40 ( .A(\SUMB[7][7] ), .Y(n130) );
  XOR2X1 U41 ( .A(n86), .B(n27), .Y(\SUMB[14][4] ) );
  XNOR2X1 U42 ( .A(\CARRYB[13][4] ), .B(\ab[14][4] ), .Y(n27) );
  XNOR2X1 U43 ( .A(n28), .B(\SUMB[12][6] ), .Y(\SUMB[13][5] ) );
  XNOR2X1 U44 ( .A(\CARRYB[12][5] ), .B(\ab[13][5] ), .Y(n28) );
  XOR2X1 U45 ( .A(n976), .B(n29), .Y(\SUMB[2][13] ) );
  XNOR2X1 U46 ( .A(\SUMB[1][14] ), .B(\ab[2][13] ), .Y(n29) );
  XNOR2X1 U47 ( .A(n30), .B(\SUMB[6][9] ), .Y(\SUMB[7][8] ) );
  XNOR2X1 U48 ( .A(\CARRYB[6][8] ), .B(\ab[7][8] ), .Y(n30) );
  XOR2X1 U49 ( .A(n158), .B(n31), .Y(n32) );
  NAND2X1 U50 ( .A(n206), .B(n1007), .Y(n31) );
  XNOR2X1 U51 ( .A(n32), .B(n271), .Y(\SUMB[2][8] ) );
  BUFX2 U52 ( .A(n883), .Y(n33) );
  XNOR2X1 U53 ( .A(\CARRYB[14][4] ), .B(n34), .Y(n676) );
  INVX8 U54 ( .A(\ab[15][4] ), .Y(n34) );
  INVX1 U55 ( .A(\SUMB[13][1] ), .Y(n35) );
  INVX1 U56 ( .A(n35), .Y(n36) );
  XOR2X1 U57 ( .A(\CARRYB[7][4] ), .B(n321), .Y(n410) );
  XOR2X1 U58 ( .A(n489), .B(n37), .Y(n267) );
  INVX8 U59 ( .A(n65), .Y(n37) );
  NAND3X1 U60 ( .A(n837), .B(n839), .C(n838), .Y(n38) );
  XOR2X1 U61 ( .A(n39), .B(n542), .Y(\SUMB[7][6] ) );
  XNOR2X1 U62 ( .A(\CARRYB[6][6] ), .B(\ab[7][6] ), .Y(n39) );
  INVX1 U63 ( .A(n1023), .Y(n40) );
  INVX2 U64 ( .A(n1022), .Y(n1023) );
  AND2X2 U65 ( .A(n810), .B(n812), .Y(n79) );
  AND2X1 U66 ( .A(n236), .B(n993), .Y(\ab[2][1] ) );
  AND2X2 U67 ( .A(n206), .B(n1007), .Y(n41) );
  XOR2X1 U68 ( .A(\SUMB[11][1] ), .B(\ab[12][0] ), .Y(n42) );
  XOR2X1 U69 ( .A(\CARRYB[11][0] ), .B(n42), .Y(\A1[10] ) );
  NAND2X1 U70 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Y(n43) );
  NAND2X1 U71 ( .A(\CARRYB[11][0] ), .B(\ab[12][0] ), .Y(n44) );
  NAND2X1 U72 ( .A(\SUMB[11][1] ), .B(\ab[12][0] ), .Y(n45) );
  NAND3X1 U73 ( .A(n44), .B(n43), .C(n45), .Y(\CARRYB[12][0] ) );
  XOR2X1 U74 ( .A(\CARRYB[3][7] ), .B(n46), .Y(n532) );
  INVX8 U75 ( .A(\ab[4][7] ), .Y(n46) );
  XOR2X1 U76 ( .A(n47), .B(n233), .Y(\SUMB[6][4] ) );
  INVX2 U77 ( .A(n47), .Y(n48) );
  INVX2 U78 ( .A(n431), .Y(n47) );
  INVX2 U79 ( .A(\SUMB[8][5] ), .Y(n253) );
  XNOR2X1 U80 ( .A(n49), .B(\SUMB[9][7] ), .Y(\SUMB[10][6] ) );
  XNOR2X1 U81 ( .A(\CARRYB[9][6] ), .B(\ab[10][6] ), .Y(n49) );
  INVX8 U82 ( .A(n52), .Y(n50) );
  INVX2 U83 ( .A(n1010), .Y(n51) );
  INVX2 U84 ( .A(B[10]), .Y(n1010) );
  INVX8 U85 ( .A(\ab[15][0] ), .Y(n52) );
  NAND3X1 U86 ( .A(n767), .B(n768), .C(n769), .Y(n53) );
  XOR2X1 U87 ( .A(n54), .B(n55), .Y(\SUMB[4][6] ) );
  XNOR2X1 U88 ( .A(\CARRYB[3][6] ), .B(\ab[4][6] ), .Y(n54) );
  INVX1 U89 ( .A(\SUMB[3][7] ), .Y(n55) );
  NAND3X1 U90 ( .A(n730), .B(n731), .C(n732), .Y(n56) );
  BUFX2 U91 ( .A(\SUMB[7][9] ), .Y(n57) );
  XOR2X1 U92 ( .A(n58), .B(n59), .Y(\SUMB[10][8] ) );
  XNOR2X1 U93 ( .A(\CARRYB[9][8] ), .B(\ab[10][8] ), .Y(n58) );
  NAND3X1 U94 ( .A(n309), .B(n308), .C(n310), .Y(n60) );
  INVX4 U95 ( .A(n996), .Y(n983) );
  INVX4 U96 ( .A(B[3]), .Y(n996) );
  INVX1 U97 ( .A(B[6]), .Y(n1002) );
  AND2X2 U98 ( .A(n439), .B(\ab[0][8] ), .Y(n61) );
  INVX4 U99 ( .A(n1004), .Y(n1005) );
  INVX4 U100 ( .A(n1010), .Y(n1011) );
  NOR2X1 U101 ( .A(n1000), .B(n40), .Y(n62) );
  AND2X2 U102 ( .A(\ab[0][3] ), .B(n964), .Y(n63) );
  XNOR2X1 U103 ( .A(\CARRYB[14][1] ), .B(n64), .Y(n561) );
  INVX8 U104 ( .A(\ab[15][1] ), .Y(n64) );
  INVX1 U105 ( .A(\CARRYB[8][6] ), .Y(n441) );
  INVX8 U106 ( .A(\ab[14][3] ), .Y(n65) );
  INVX2 U107 ( .A(\ab[10][5] ), .Y(n157) );
  INVX2 U108 ( .A(\ab[11][4] ), .Y(n301) );
  INVX2 U109 ( .A(\ab[4][9] ), .Y(n401) );
  INVX2 U110 ( .A(\ab[12][3] ), .Y(n149) );
  INVX2 U111 ( .A(\ab[6][7] ), .Y(n205) );
  INVX2 U112 ( .A(\ab[5][7] ), .Y(n261) );
  INVX2 U113 ( .A(\ab[7][7] ), .Y(n440) );
  INVX2 U114 ( .A(\ab[12][6] ), .Y(n244) );
  INVX2 U115 ( .A(\ab[7][10] ), .Y(n248) );
  INVX2 U116 ( .A(\ab[11][5] ), .Y(n298) );
  INVX2 U117 ( .A(\ab[10][4] ), .Y(n163) );
  INVX2 U118 ( .A(\ab[13][2] ), .Y(n251) );
  INVX2 U119 ( .A(\ab[14][6] ), .Y(n186) );
  INVX2 U120 ( .A(\ab[6][9] ), .Y(n138) );
  INVX2 U121 ( .A(\ab[6][8] ), .Y(n175) );
  INVX2 U122 ( .A(\ab[4][5] ), .Y(n182) );
  INVX2 U123 ( .A(\ab[7][5] ), .Y(n503) );
  INVX2 U124 ( .A(\ab[9][5] ), .Y(n224) );
  INVX2 U125 ( .A(\ab[8][3] ), .Y(n755) );
  INVX2 U126 ( .A(\ab[8][4] ), .Y(n321) );
  INVX2 U127 ( .A(\ab[9][9] ), .Y(n189) );
  INVX4 U128 ( .A(n1002), .Y(n1003) );
  INVX2 U129 ( .A(\ab[14][1] ), .Y(n530) );
  INVX2 U130 ( .A(n318), .Y(n317) );
  INVX2 U131 ( .A(\ab[13][8] ), .Y(n324) );
  AND2X1 U132 ( .A(\SUMB[15][8] ), .B(\CARRYB[15][7] ), .Y(n66) );
  AND2X2 U133 ( .A(\SUMB[15][9] ), .B(\CARRYB[15][8] ), .Y(n67) );
  AND2X2 U134 ( .A(\SUMB[15][10] ), .B(\CARRYB[15][9] ), .Y(n68) );
  AND2X2 U135 ( .A(\SUMB[15][11] ), .B(\CARRYB[15][10] ), .Y(n69) );
  AND2X2 U136 ( .A(\SUMB[15][12] ), .B(\CARRYB[15][11] ), .Y(n70) );
  AND2X2 U137 ( .A(\SUMB[15][13] ), .B(\CARRYB[15][12] ), .Y(n71) );
  AND2X2 U138 ( .A(\SUMB[15][14] ), .B(\CARRYB[15][13] ), .Y(n72) );
  AND2X2 U139 ( .A(\SUMB[15][15] ), .B(\CARRYB[15][14] ), .Y(n73) );
  AND2X2 U140 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n74) );
  AND2X2 U141 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Y(n75) );
  XOR2X1 U142 ( .A(\SUMB[10][8] ), .B(n586), .Y(n76) );
  AND2X2 U143 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(n77) );
  AND2X2 U144 ( .A(n527), .B(n529), .Y(n78) );
  AND2X2 U145 ( .A(\SUMB[15][7] ), .B(\CARRYB[15][6] ), .Y(n80) );
  XNOR2X1 U146 ( .A(n81), .B(\SUMB[2][10] ), .Y(\SUMB[3][9] ) );
  XNOR2X1 U147 ( .A(\CARRYB[2][9] ), .B(\ab[3][9] ), .Y(n81) );
  AND2X2 U148 ( .A(n236), .B(n1013), .Y(n82) );
  XNOR2X1 U149 ( .A(\ab[0][10] ), .B(n83), .Y(\SUMB[1][9] ) );
  NAND2X1 U150 ( .A(B[9]), .B(n322), .Y(n83) );
  NAND3X1 U151 ( .A(n887), .B(n888), .C(n889), .Y(n84) );
  NAND3X1 U152 ( .A(n404), .B(n403), .C(n405), .Y(n85) );
  INVX2 U153 ( .A(\CARRYB[15][5] ), .Y(n318) );
  INVX1 U154 ( .A(\SUMB[13][5] ), .Y(n86) );
  NAND3X1 U155 ( .A(n714), .B(n715), .C(n716), .Y(n87) );
  BUFX2 U156 ( .A(n638), .Y(n88) );
  BUFX2 U157 ( .A(\SUMB[9][1] ), .Y(n89) );
  XOR2X1 U158 ( .A(n90), .B(n272), .Y(\SUMB[6][7] ) );
  XOR2X1 U159 ( .A(\SUMB[5][8] ), .B(n205), .Y(n90) );
  NAND3X1 U160 ( .A(n679), .B(n678), .C(n677), .Y(\CARRYB[15][4] ) );
  XOR2X1 U161 ( .A(n91), .B(n57), .Y(\SUMB[8][8] ) );
  XOR2X1 U162 ( .A(\CARRYB[7][8] ), .B(\ab[8][8] ), .Y(n91) );
  BUFX2 U163 ( .A(\CARRYB[7][2] ), .Y(n92) );
  XOR2X1 U164 ( .A(n311), .B(n312), .Y(n93) );
  INVX2 U165 ( .A(\SUMB[10][5] ), .Y(n311) );
  BUFX2 U166 ( .A(\CARRYB[3][10] ), .Y(n94) );
  XOR2X1 U167 ( .A(n152), .B(n128), .Y(n95) );
  BUFX2 U168 ( .A(\CARRYB[3][5] ), .Y(n96) );
  XOR2X1 U169 ( .A(n172), .B(n215), .Y(n97) );
  NAND3X1 U170 ( .A(n675), .B(n673), .C(n674), .Y(n98) );
  NAND3X1 U171 ( .A(n778), .B(n779), .C(n780), .Y(n99) );
  XOR2X1 U172 ( .A(n410), .B(n534), .Y(n100) );
  INVX2 U173 ( .A(\SUMB[7][5] ), .Y(n534) );
  XOR2X1 U174 ( .A(\CARRYB[9][3] ), .B(\ab[10][3] ), .Y(n449) );
  AND2X2 U175 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(n737) );
  XOR2X1 U176 ( .A(\CARRYB[5][13] ), .B(\ab[6][13] ), .Y(n101) );
  XOR2X1 U177 ( .A(\SUMB[5][14] ), .B(n101), .Y(\SUMB[6][13] ) );
  NAND2X1 U178 ( .A(\SUMB[5][14] ), .B(\CARRYB[5][13] ), .Y(n102) );
  NAND2X1 U179 ( .A(\SUMB[5][14] ), .B(\ab[6][13] ), .Y(n103) );
  NAND2X1 U180 ( .A(\CARRYB[5][13] ), .B(\ab[6][13] ), .Y(n104) );
  NAND3X1 U181 ( .A(n103), .B(n102), .C(n104), .Y(\CARRYB[6][13] ) );
  XOR2X1 U182 ( .A(\ab[5][14] ), .B(\ab[4][15] ), .Y(n105) );
  XOR2X1 U183 ( .A(\CARRYB[4][14] ), .B(n105), .Y(\SUMB[5][14] ) );
  NAND2X1 U184 ( .A(\CARRYB[4][14] ), .B(\ab[5][14] ), .Y(n106) );
  NAND2X1 U185 ( .A(\CARRYB[4][14] ), .B(\ab[4][15] ), .Y(n107) );
  NAND2X1 U186 ( .A(\ab[5][14] ), .B(\ab[4][15] ), .Y(n108) );
  NAND3X1 U187 ( .A(n107), .B(n106), .C(n108), .Y(\CARRYB[5][14] ) );
  XOR2X1 U188 ( .A(\CARRYB[13][8] ), .B(\ab[14][8] ), .Y(n109) );
  XOR2X1 U189 ( .A(\SUMB[13][9] ), .B(n109), .Y(\SUMB[14][8] ) );
  NAND2X1 U190 ( .A(\SUMB[13][9] ), .B(\CARRYB[13][8] ), .Y(n110) );
  NAND2X1 U191 ( .A(\SUMB[13][9] ), .B(\ab[14][8] ), .Y(n111) );
  NAND2X1 U192 ( .A(\CARRYB[13][8] ), .B(\ab[14][8] ), .Y(n112) );
  NAND3X1 U193 ( .A(n111), .B(n110), .C(n112), .Y(\CARRYB[14][8] ) );
  XOR2X1 U194 ( .A(\CARRYB[10][10] ), .B(\ab[11][10] ), .Y(n113) );
  XOR2X1 U195 ( .A(\SUMB[10][11] ), .B(n113), .Y(\SUMB[11][10] ) );
  NAND2X1 U196 ( .A(\SUMB[10][11] ), .B(\CARRYB[10][10] ), .Y(n114) );
  NAND2X1 U197 ( .A(\SUMB[10][11] ), .B(\ab[11][10] ), .Y(n115) );
  NAND2X1 U198 ( .A(\CARRYB[10][10] ), .B(\ab[11][10] ), .Y(n116) );
  NAND3X1 U199 ( .A(n115), .B(n114), .C(n116), .Y(\CARRYB[11][10] ) );
  BUFX2 U200 ( .A(\SUMB[6][12] ), .Y(n117) );
  XNOR2X1 U201 ( .A(n118), .B(\SUMB[5][13] ), .Y(\SUMB[6][12] ) );
  XOR2X1 U202 ( .A(n711), .B(\ab[6][12] ), .Y(n118) );
  XOR2X1 U203 ( .A(\SUMB[15][5] ), .B(\CARRYB[15][4] ), .Y(\A1[18] ) );
  BUFX2 U204 ( .A(n748), .Y(n119) );
  BUFX2 U205 ( .A(n794), .Y(n120) );
  BUFX2 U206 ( .A(\SUMB[4][5] ), .Y(n121) );
  NAND3X1 U207 ( .A(n666), .B(n664), .C(n665), .Y(n122) );
  XOR2X1 U208 ( .A(\CARRYB[10][7] ), .B(\ab[11][7] ), .Y(n586) );
  XOR2X1 U209 ( .A(\CARRYB[12][6] ), .B(\ab[13][6] ), .Y(n424) );
  BUFX2 U210 ( .A(n698), .Y(n123) );
  NAND3X1 U211 ( .A(n587), .B(n588), .C(n589), .Y(n124) );
  XNOR2X1 U212 ( .A(n125), .B(\SUMB[12][8] ), .Y(\SUMB[13][7] ) );
  XNOR2X1 U213 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .Y(n125) );
  NAND3X1 U214 ( .A(n667), .B(n668), .C(n669), .Y(n126) );
  XOR2X1 U215 ( .A(\SUMB[8][9] ), .B(n127), .Y(\SUMB[9][8] ) );
  XOR2X1 U216 ( .A(\CARRYB[8][8] ), .B(\ab[9][8] ), .Y(n127) );
  XOR2X1 U217 ( .A(n152), .B(n128), .Y(\SUMB[5][11] ) );
  XOR2X1 U218 ( .A(\CARRYB[4][11] ), .B(\ab[5][11] ), .Y(n128) );
  XOR2X1 U219 ( .A(n129), .B(n130), .Y(\SUMB[8][6] ) );
  XNOR2X1 U220 ( .A(n147), .B(\ab[8][6] ), .Y(n129) );
  INVX1 U221 ( .A(n1007), .Y(n131) );
  INVX4 U222 ( .A(n131), .Y(n132) );
  INVX4 U223 ( .A(n1006), .Y(n1007) );
  INVX2 U224 ( .A(B[8]), .Y(n1006) );
  XOR2X1 U225 ( .A(\SUMB[11][2] ), .B(\ab[12][1] ), .Y(n169) );
  XNOR2X1 U226 ( .A(n133), .B(n100), .Y(\SUMB[9][3] ) );
  XNOR2X1 U227 ( .A(\CARRYB[8][3] ), .B(\ab[9][3] ), .Y(n133) );
  XNOR2X1 U228 ( .A(n134), .B(n135), .Y(\SUMB[11][2] ) );
  XOR2X1 U229 ( .A(\CARRYB[10][2] ), .B(\ab[11][2] ), .Y(n134) );
  XOR2X1 U230 ( .A(n449), .B(n377), .Y(n135) );
  INVX2 U231 ( .A(\SUMB[6][7] ), .Y(n542) );
  XNOR2X1 U232 ( .A(n136), .B(\SUMB[12][3] ), .Y(\SUMB[13][2] ) );
  XOR2X1 U233 ( .A(\CARRYB[12][2] ), .B(n251), .Y(n136) );
  XNOR2X1 U234 ( .A(\ab[1][11] ), .B(n137), .Y(\SUMB[1][11] ) );
  NAND2X1 U235 ( .A(n266), .B(n1015), .Y(n137) );
  XNOR2X1 U236 ( .A(n336), .B(n138), .Y(n726) );
  INVX1 U237 ( .A(\SUMB[5][5] ), .Y(n431) );
  INVX1 U238 ( .A(n974), .Y(\CARRYB[1][9] ) );
  XNOR2X1 U239 ( .A(n725), .B(n139), .Y(\SUMB[5][10] ) );
  INVX2 U240 ( .A(\SUMB[4][11] ), .Y(n139) );
  AND2X1 U241 ( .A(\SUMB[15][4] ), .B(\CARRYB[15][3] ), .Y(n967) );
  XOR2X1 U242 ( .A(\SUMB[1][5] ), .B(\ab[2][4] ), .Y(n140) );
  XOR2X1 U243 ( .A(n965), .B(n140), .Y(\SUMB[2][4] ) );
  NAND2X1 U244 ( .A(n965), .B(\SUMB[1][5] ), .Y(n141) );
  NAND2X1 U245 ( .A(n965), .B(\ab[2][4] ), .Y(n142) );
  NAND2X1 U246 ( .A(\SUMB[1][5] ), .B(\ab[2][4] ), .Y(n143) );
  NAND3X1 U247 ( .A(n142), .B(n141), .C(n143), .Y(\CARRYB[2][4] ) );
  BUFX2 U248 ( .A(\CARRYB[12][0] ), .Y(n144) );
  NAND3X1 U249 ( .A(n870), .B(n869), .C(n871), .Y(n145) );
  BUFX2 U250 ( .A(\SUMB[9][6] ), .Y(n146) );
  NAND3X1 U251 ( .A(n944), .B(n943), .C(n942), .Y(n147) );
  INVX1 U252 ( .A(\SUMB[5][10] ), .Y(n300) );
  AND2X2 U253 ( .A(n266), .B(n1015), .Y(n148) );
  XOR2X1 U254 ( .A(\CARRYB[11][3] ), .B(n149), .Y(n195) );
  INVX2 U255 ( .A(n1022), .Y(n235) );
  INVX2 U256 ( .A(n1022), .Y(n236) );
  INVX1 U257 ( .A(\SUMB[1][14] ), .Y(n150) );
  INVX1 U258 ( .A(n150), .Y(n151) );
  BUFX2 U259 ( .A(\SUMB[4][12] ), .Y(n152) );
  XOR2X1 U260 ( .A(\SUMB[8][11] ), .B(\ab[9][10] ), .Y(n153) );
  XOR2X1 U261 ( .A(n153), .B(\CARRYB[8][10] ), .Y(\SUMB[9][10] ) );
  NAND2X1 U262 ( .A(\CARRYB[8][10] ), .B(\SUMB[8][11] ), .Y(n154) );
  NAND2X1 U263 ( .A(\CARRYB[8][10] ), .B(\ab[9][10] ), .Y(n155) );
  NAND2X1 U264 ( .A(\SUMB[8][11] ), .B(\ab[9][10] ), .Y(n156) );
  NAND3X1 U265 ( .A(n155), .B(n154), .C(n156), .Y(\CARRYB[9][10] ) );
  INVX1 U266 ( .A(n472), .Y(n473) );
  INVX2 U267 ( .A(\SUMB[1][9] ), .Y(n271) );
  NAND2X1 U268 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(n158) );
  XOR2X1 U269 ( .A(n159), .B(n160), .Y(\SUMB[6][1] ) );
  XNOR2X1 U270 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .Y(n159) );
  INVX1 U271 ( .A(\SUMB[5][2] ), .Y(n160) );
  XNOR2X1 U272 ( .A(n791), .B(n161), .Y(\SUMB[7][9] ) );
  INVX2 U273 ( .A(\SUMB[6][10] ), .Y(n161) );
  AND2X2 U274 ( .A(\CARRYB[15][1] ), .B(\SUMB[15][2] ), .Y(n971) );
  BUFX2 U275 ( .A(n835), .Y(n162) );
  XOR2X1 U276 ( .A(\CARRYB[9][4] ), .B(n163), .Y(n376) );
  BUFX2 U277 ( .A(\SUMB[8][1] ), .Y(n164) );
  XOR2X1 U278 ( .A(\CARRYB[10][1] ), .B(\ab[11][1] ), .Y(n165) );
  XOR2X1 U279 ( .A(n165), .B(\SUMB[10][2] ), .Y(\SUMB[11][1] ) );
  XNOR2X1 U280 ( .A(n166), .B(\SUMB[14][3] ), .Y(\SUMB[15][2] ) );
  XNOR2X1 U281 ( .A(\CARRYB[14][2] ), .B(\ab[15][2] ), .Y(n166) );
  XOR2X1 U282 ( .A(n167), .B(\SUMB[13][7] ), .Y(\SUMB[14][6] ) );
  XNOR2X1 U283 ( .A(\CARRYB[13][6] ), .B(n186), .Y(n167) );
  XNOR2X1 U284 ( .A(n168), .B(n171), .Y(\SUMB[7][5] ) );
  XOR2X1 U285 ( .A(\SUMB[6][6] ), .B(n503), .Y(n168) );
  XNOR2X1 U286 ( .A(n169), .B(n170), .Y(\SUMB[12][1] ) );
  INVX1 U287 ( .A(\CARRYB[11][1] ), .Y(n170) );
  BUFX2 U288 ( .A(\CARRYB[6][5] ), .Y(n171) );
  XOR2X1 U289 ( .A(n172), .B(n215), .Y(\SUMB[2][7] ) );
  XNOR2X1 U290 ( .A(n435), .B(n314), .Y(n172) );
  INVX1 U291 ( .A(\CARRYB[2][8] ), .Y(n436) );
  NAND3X1 U292 ( .A(n803), .B(n802), .C(n801), .Y(n173) );
  NAND3X1 U293 ( .A(n885), .B(n884), .C(n886), .Y(n174) );
  XNOR2X1 U294 ( .A(n176), .B(\SUMB[7][8] ), .Y(\SUMB[8][7] ) );
  XNOR2X1 U295 ( .A(\CARRYB[7][7] ), .B(\ab[8][7] ), .Y(n176) );
  XNOR2X1 U296 ( .A(n177), .B(n223), .Y(\SUMB[3][10] ) );
  XNOR2X1 U297 ( .A(\CARRYB[2][10] ), .B(\ab[3][10] ), .Y(n177) );
  INVX2 U298 ( .A(n998), .Y(n984) );
  INVX4 U299 ( .A(n986), .Y(n514) );
  XOR2X1 U300 ( .A(n178), .B(\CARRYB[5][2] ), .Y(\SUMB[6][2] ) );
  XOR2X1 U301 ( .A(\SUMB[5][3] ), .B(\ab[6][2] ), .Y(n178) );
  NAND3X1 U302 ( .A(n257), .B(n258), .C(n259), .Y(n179) );
  NAND3X1 U303 ( .A(n383), .B(n382), .C(n384), .Y(n180) );
  AND2X2 U304 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n181) );
  AND2X2 U305 ( .A(B[6]), .B(n987), .Y(n524) );
  XOR2X1 U306 ( .A(\SUMB[3][6] ), .B(n182), .Y(n234) );
  XOR2X1 U307 ( .A(n183), .B(n97), .Y(\SUMB[3][6] ) );
  XNOR2X1 U308 ( .A(n847), .B(\ab[3][6] ), .Y(n183) );
  XOR2X1 U309 ( .A(\CARRYB[7][3] ), .B(n755), .Y(n216) );
  AND2X2 U310 ( .A(B[9]), .B(n322), .Y(n184) );
  BUFX2 U311 ( .A(\CARRYB[4][3] ), .Y(n185) );
  BUFX2 U312 ( .A(n894), .Y(n187) );
  INVX2 U313 ( .A(\SUMB[8][3] ), .Y(n608) );
  XOR2X1 U314 ( .A(n448), .B(n188), .Y(\SUMB[8][5] ) );
  INVX2 U315 ( .A(\SUMB[7][6] ), .Y(n188) );
  XOR2X1 U316 ( .A(n189), .B(n220), .Y(n194) );
  INVX1 U317 ( .A(n220), .Y(n221) );
  NAND3X1 U318 ( .A(n955), .B(n954), .C(n956), .Y(n190) );
  XNOR2X1 U319 ( .A(n191), .B(n192), .Y(\SUMB[7][3] ) );
  XOR2X1 U320 ( .A(n413), .B(\ab[7][3] ), .Y(n191) );
  XOR2X1 U321 ( .A(n233), .B(n48), .Y(n192) );
  NAND3X1 U322 ( .A(n479), .B(n478), .C(n480), .Y(n193) );
  INVX1 U323 ( .A(\CARRYB[6][2] ), .Y(n960) );
  XOR2X1 U324 ( .A(n194), .B(\SUMB[8][10] ), .Y(\SUMB[9][9] ) );
  XNOR2X1 U325 ( .A(n195), .B(n93), .Y(\SUMB[12][3] ) );
  BUFX2 U326 ( .A(\SUMB[3][5] ), .Y(n196) );
  NAND3X1 U327 ( .A(n958), .B(n959), .C(n957), .Y(n197) );
  XOR2X1 U328 ( .A(\SUMB[3][11] ), .B(\ab[4][10] ), .Y(n198) );
  XOR2X1 U329 ( .A(n94), .B(n198), .Y(\SUMB[4][10] ) );
  NAND2X1 U330 ( .A(\SUMB[3][11] ), .B(\CARRYB[3][10] ), .Y(n199) );
  NAND2X1 U331 ( .A(\CARRYB[3][10] ), .B(\ab[4][10] ), .Y(n200) );
  NAND2X1 U332 ( .A(\SUMB[3][11] ), .B(\ab[4][10] ), .Y(n201) );
  NAND3X1 U333 ( .A(n200), .B(n199), .C(n201), .Y(\CARRYB[4][10] ) );
  NAND3X1 U334 ( .A(n624), .B(n625), .C(n626), .Y(n202) );
  NAND3X1 U335 ( .A(n764), .B(n13), .C(n766), .Y(n203) );
  NAND3X1 U336 ( .A(n834), .B(n836), .C(n162), .Y(n204) );
  INVX2 U337 ( .A(n1022), .Y(n206) );
  XOR2X1 U338 ( .A(n207), .B(n208), .Y(\SUMB[7][4] ) );
  XNOR2X1 U339 ( .A(n122), .B(\ab[7][4] ), .Y(n207) );
  INVX2 U340 ( .A(\SUMB[6][5] ), .Y(n208) );
  XOR2X1 U341 ( .A(\SUMB[3][14] ), .B(\ab[4][13] ), .Y(n209) );
  XOR2X1 U342 ( .A(\CARRYB[3][13] ), .B(n209), .Y(\SUMB[4][13] ) );
  NAND2X1 U343 ( .A(\CARRYB[3][13] ), .B(\SUMB[3][14] ), .Y(n210) );
  NAND2X1 U344 ( .A(\CARRYB[3][13] ), .B(\ab[4][13] ), .Y(n211) );
  NAND2X1 U345 ( .A(\SUMB[3][14] ), .B(\ab[4][13] ), .Y(n212) );
  NAND3X1 U346 ( .A(n211), .B(n210), .C(n212), .Y(\CARRYB[4][13] ) );
  NAND3X1 U347 ( .A(n391), .B(n390), .C(n392), .Y(n213) );
  INVX1 U348 ( .A(n847), .Y(n848) );
  INVX1 U349 ( .A(\SUMB[1][12] ), .Y(n297) );
  XOR2X1 U350 ( .A(n219), .B(n269), .Y(n214) );
  BUFX2 U351 ( .A(\SUMB[1][8] ), .Y(n215) );
  XOR2X1 U352 ( .A(n216), .B(n375), .Y(\SUMB[8][3] ) );
  XNOR2X1 U353 ( .A(n519), .B(n217), .Y(\SUMB[2][6] ) );
  INVX1 U354 ( .A(\SUMB[1][7] ), .Y(n217) );
  NAND2X1 U355 ( .A(n1025), .B(n1007), .Y(n218) );
  INVX2 U356 ( .A(n218), .Y(\ab[3][8] ) );
  XOR2X1 U357 ( .A(n269), .B(n219), .Y(\SUMB[3][12] ) );
  XNOR2X1 U358 ( .A(\CARRYB[2][12] ), .B(\ab[3][12] ), .Y(n219) );
  INVX2 U359 ( .A(\CARRYB[8][9] ), .Y(n220) );
  AND2X2 U360 ( .A(n148), .B(\ab[1][11] ), .Y(n222) );
  XOR2X1 U361 ( .A(n615), .B(\SUMB[2][9] ), .Y(\SUMB[3][8] ) );
  BUFX2 U362 ( .A(n895), .Y(n225) );
  XOR2X1 U363 ( .A(n226), .B(\SUMB[6][8] ), .Y(\SUMB[7][7] ) );
  XNOR2X1 U364 ( .A(\CARRYB[6][7] ), .B(n440), .Y(n226) );
  INVX1 U365 ( .A(\SUMB[15][5] ), .Y(n227) );
  INVX1 U366 ( .A(n227), .Y(n228) );
  XNOR2X1 U367 ( .A(n229), .B(n214), .Y(\SUMB[4][11] ) );
  XNOR2X1 U368 ( .A(\CARRYB[3][11] ), .B(\ab[4][11] ), .Y(n229) );
  INVX1 U369 ( .A(n445), .Y(n230) );
  NAND3X1 U370 ( .A(n576), .B(n578), .C(n577), .Y(n231) );
  XNOR2X1 U371 ( .A(n232), .B(\SUMB[2][12] ), .Y(\SUMB[3][11] ) );
  XNOR2X1 U372 ( .A(\CARRYB[2][11] ), .B(\ab[3][11] ), .Y(n232) );
  XOR2X1 U373 ( .A(n975), .B(\ab[2][12] ), .Y(n252) );
  INVX1 U374 ( .A(n975), .Y(\CARRYB[1][12] ) );
  XOR2X1 U375 ( .A(\CARRYB[5][4] ), .B(\ab[6][4] ), .Y(n233) );
  XNOR2X1 U376 ( .A(n234), .B(n96), .Y(\SUMB[4][5] ) );
  BUFX2 U377 ( .A(n601), .Y(n237) );
  NAND3X1 U378 ( .A(n872), .B(n873), .C(n874), .Y(n238) );
  INVX1 U379 ( .A(n1006), .Y(n239) );
  BUFX2 U380 ( .A(\CARRYB[10][0] ), .Y(n240) );
  BUFX2 U381 ( .A(n663), .Y(n241) );
  INVX1 U382 ( .A(n486), .Y(n242) );
  INVX1 U383 ( .A(n242), .Y(n243) );
  NAND3X1 U384 ( .A(n822), .B(n823), .C(n824), .Y(n245) );
  NAND3X1 U385 ( .A(n828), .B(n830), .C(n829), .Y(n246) );
  XOR2X1 U386 ( .A(n411), .B(n412), .Y(n247) );
  AND2X2 U387 ( .A(ZB), .B(n1020), .Y(\ab[0][15] ) );
  XOR2X1 U388 ( .A(\CARRYB[6][10] ), .B(n248), .Y(n750) );
  INVX2 U389 ( .A(\SUMB[9][8] ), .Y(n736) );
  XOR2X1 U390 ( .A(n249), .B(n250), .Y(\SUMB[6][11] ) );
  XNOR2X1 U391 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .Y(n249) );
  INVX2 U392 ( .A(\SUMB[5][12] ), .Y(n250) );
  XNOR2X1 U393 ( .A(n252), .B(\SUMB[1][13] ), .Y(\SUMB[2][12] ) );
  NAND2X1 U394 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .Y(n254) );
  NAND2X1 U395 ( .A(\SUMB[7][7] ), .B(\ab[8][6] ), .Y(n255) );
  NAND2X1 U396 ( .A(\CARRYB[7][6] ), .B(\SUMB[7][7] ), .Y(n256) );
  NAND3X1 U397 ( .A(n254), .B(n255), .C(n256), .Y(\CARRYB[8][6] ) );
  NAND2X1 U398 ( .A(n204), .B(\ab[9][5] ), .Y(n257) );
  NAND2X1 U399 ( .A(\SUMB[8][6] ), .B(\ab[9][5] ), .Y(n258) );
  NAND2X1 U400 ( .A(n204), .B(\SUMB[8][6] ), .Y(n259) );
  NAND3X1 U401 ( .A(n257), .B(n258), .C(n259), .Y(\CARRYB[9][5] ) );
  NAND3X1 U402 ( .A(n641), .B(n642), .C(n643), .Y(n260) );
  XOR2X1 U403 ( .A(\CARRYB[4][7] ), .B(n261), .Y(n543) );
  NAND2X1 U404 ( .A(\ab[6][5] ), .B(n263), .Y(n264) );
  NAND2X1 U405 ( .A(n262), .B(n245), .Y(n265) );
  NAND2X1 U406 ( .A(n264), .B(n265), .Y(n700) );
  INVX1 U407 ( .A(\ab[6][5] ), .Y(n262) );
  INVX1 U408 ( .A(\CARRYB[5][5] ), .Y(n263) );
  INVX4 U409 ( .A(B[12]), .Y(n1014) );
  INVX2 U410 ( .A(\CARRYB[5][7] ), .Y(n272) );
  BUFX4 U411 ( .A(A[0]), .Y(n266) );
  INVX2 U412 ( .A(A[0]), .Y(n1020) );
  XNOR2X1 U413 ( .A(n267), .B(n268), .Y(\SUMB[14][3] ) );
  INVX2 U414 ( .A(\SUMB[13][4] ), .Y(n268) );
  INVX2 U415 ( .A(\SUMB[2][13] ), .Y(n269) );
  NAND3X1 U416 ( .A(n843), .B(n845), .C(n844), .Y(n270) );
  XNOR2X1 U417 ( .A(n273), .B(n274), .Y(\SUMB[13][3] ) );
  XOR2X1 U418 ( .A(\CARRYB[12][3] ), .B(\ab[13][3] ), .Y(n273) );
  XNOR2X1 U419 ( .A(n339), .B(n414), .Y(n274) );
  INVX1 U420 ( .A(\SUMB[7][2] ), .Y(n373) );
  NAND3X1 U421 ( .A(n661), .B(n662), .C(n241), .Y(n275) );
  NAND3X1 U422 ( .A(n717), .B(n718), .C(n719), .Y(n276) );
  NAND3X1 U423 ( .A(n602), .B(n603), .C(n604), .Y(n277) );
  NAND3X1 U424 ( .A(n878), .B(n879), .C(n880), .Y(n278) );
  NAND3X1 U425 ( .A(n537), .B(n536), .C(n538), .Y(n279) );
  BUFX2 U426 ( .A(n793), .Y(n280) );
  XNOR2X1 U427 ( .A(n281), .B(\SUMB[11][8] ), .Y(\SUMB[12][7] ) );
  XNOR2X1 U428 ( .A(\CARRYB[11][7] ), .B(\ab[12][7] ), .Y(n281) );
  XOR2X1 U429 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .Y(n282) );
  XOR2X1 U430 ( .A(n282), .B(\SUMB[13][8] ), .Y(\SUMB[14][7] ) );
  XOR2X1 U431 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .Y(n283) );
  XOR2X1 U432 ( .A(n283), .B(\SUMB[14][7] ), .Y(\SUMB[15][6] ) );
  NAND2X1 U433 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .Y(n284) );
  NAND2X1 U434 ( .A(\ab[14][7] ), .B(\SUMB[13][8] ), .Y(n285) );
  NAND2X1 U435 ( .A(\CARRYB[13][7] ), .B(\SUMB[13][8] ), .Y(n286) );
  NAND3X1 U436 ( .A(n284), .B(n285), .C(n286), .Y(\CARRYB[14][7] ) );
  NAND2X1 U437 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .Y(n287) );
  NAND2X1 U438 ( .A(\ab[15][6] ), .B(\SUMB[14][7] ), .Y(n288) );
  NAND2X1 U439 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Y(n289) );
  NAND3X1 U440 ( .A(n287), .B(n288), .C(n289), .Y(\CARRYB[15][6] ) );
  XOR2X1 U441 ( .A(\CARRYB[11][8] ), .B(\ab[12][8] ), .Y(n290) );
  XOR2X1 U442 ( .A(\SUMB[11][9] ), .B(n290), .Y(\SUMB[12][8] ) );
  NAND2X1 U443 ( .A(\SUMB[11][9] ), .B(n213), .Y(n291) );
  NAND2X1 U444 ( .A(\SUMB[11][9] ), .B(\ab[12][8] ), .Y(n292) );
  NAND2X1 U445 ( .A(n213), .B(\ab[12][8] ), .Y(n293) );
  NAND3X1 U446 ( .A(n292), .B(n291), .C(n293), .Y(\CARRYB[12][8] ) );
  BUFX2 U447 ( .A(\CARRYB[4][12] ), .Y(n294) );
  NAND3X1 U448 ( .A(n684), .B(n685), .C(n686), .Y(n295) );
  INVX2 U449 ( .A(\SUMB[1][10] ), .Y(n337) );
  XOR2X1 U450 ( .A(\CARRYB[13][5] ), .B(\ab[14][5] ), .Y(n332) );
  XNOR2X1 U451 ( .A(n296), .B(n736), .Y(\SUMB[10][7] ) );
  XOR2X1 U452 ( .A(\CARRYB[9][7] ), .B(\ab[10][7] ), .Y(n296) );
  XNOR2X1 U453 ( .A(\CARRYB[10][5] ), .B(n298), .Y(n598) );
  NAND3X1 U454 ( .A(n893), .B(n225), .C(n187), .Y(n299) );
  XNOR2X1 U455 ( .A(n726), .B(n300), .Y(\SUMB[6][9] ) );
  INVX8 U456 ( .A(ZB), .Y(n1049) );
  XOR2X1 U457 ( .A(\CARRYB[10][4] ), .B(n301), .Y(n312) );
  NAND3X1 U458 ( .A(n825), .B(n826), .C(n827), .Y(n302) );
  NAND3X1 U459 ( .A(n832), .B(n831), .C(n833), .Y(n303) );
  XOR2X1 U460 ( .A(\SUMB[4][13] ), .B(\ab[5][12] ), .Y(n304) );
  XOR2X1 U461 ( .A(n304), .B(n294), .Y(\SUMB[5][12] ) );
  NAND2X1 U462 ( .A(\CARRYB[4][12] ), .B(\SUMB[4][13] ), .Y(n305) );
  NAND2X1 U463 ( .A(\CARRYB[4][12] ), .B(\ab[5][12] ), .Y(n306) );
  NAND2X1 U464 ( .A(\SUMB[4][13] ), .B(\ab[5][12] ), .Y(n307) );
  NAND3X1 U465 ( .A(n307), .B(n305), .C(n306), .Y(\CARRYB[5][12] ) );
  NAND2X1 U466 ( .A(\SUMB[1][14] ), .B(\CARRYB[1][13] ), .Y(n308) );
  NAND2X1 U467 ( .A(\CARRYB[1][13] ), .B(\ab[2][13] ), .Y(n309) );
  NAND2X1 U468 ( .A(n151), .B(\ab[2][13] ), .Y(n310) );
  NAND3X1 U469 ( .A(n309), .B(n308), .C(n310), .Y(\CARRYB[2][13] ) );
  NAND3X1 U470 ( .A(n804), .B(n805), .C(n806), .Y(n313) );
  INVX2 U471 ( .A(n1021), .Y(n846) );
  NAND2X1 U472 ( .A(\ab[0][8] ), .B(n439), .Y(n314) );
  BUFX2 U473 ( .A(\SUMB[15][0] ), .Y(n315) );
  NAND3X1 U474 ( .A(n500), .B(n501), .C(n502), .Y(n316) );
  XOR2X1 U475 ( .A(\SUMB[15][6] ), .B(n317), .Y(\A1[19] ) );
  XNOR2X1 U476 ( .A(n319), .B(\SUMB[7][12] ), .Y(\SUMB[8][11] ) );
  XNOR2X1 U477 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .Y(n319) );
  XOR2X1 U478 ( .A(n474), .B(n320), .Y(\SUMB[13][1] ) );
  BUFX2 U479 ( .A(A[1]), .Y(n322) );
  INVX1 U480 ( .A(A[1]), .Y(n1021) );
  XNOR2X1 U481 ( .A(\ab[7][12] ), .B(n712), .Y(n680) );
  INVX1 U482 ( .A(n712), .Y(n713) );
  INVX1 U483 ( .A(n441), .Y(n442) );
  XNOR2X1 U484 ( .A(n323), .B(n77), .Y(\SUMB[2][10] ) );
  XNOR2X1 U485 ( .A(\SUMB[1][11] ), .B(\ab[2][10] ), .Y(n323) );
  XNOR2X1 U486 ( .A(n324), .B(\CARRYB[12][8] ), .Y(n457) );
  XNOR2X1 U487 ( .A(n325), .B(n326), .Y(\SUMB[12][2] ) );
  XOR2X1 U488 ( .A(\CARRYB[11][2] ), .B(\ab[12][2] ), .Y(n325) );
  XNOR2X1 U489 ( .A(n10), .B(n374), .Y(n326) );
  XNOR2X1 U490 ( .A(n327), .B(\SUMB[2][14] ), .Y(\SUMB[3][13] ) );
  XNOR2X1 U491 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .Y(n327) );
  NAND3X1 U492 ( .A(n599), .B(n600), .C(n237), .Y(n328) );
  NAND3X1 U493 ( .A(n896), .B(n897), .C(n24), .Y(n329) );
  NAND3X1 U494 ( .A(n658), .B(n660), .C(n659), .Y(n330) );
  XOR2X1 U495 ( .A(n763), .B(n374), .Y(n331) );
  XOR2X1 U496 ( .A(n332), .B(\SUMB[13][6] ), .Y(\SUMB[14][5] ) );
  NAND2X1 U497 ( .A(\SUMB[13][6] ), .B(n99), .Y(n333) );
  NAND2X1 U498 ( .A(\SUMB[13][6] ), .B(\ab[14][5] ), .Y(n334) );
  NAND2X1 U499 ( .A(n99), .B(\ab[14][5] ), .Y(n335) );
  NAND3X1 U500 ( .A(n334), .B(n333), .C(n335), .Y(\CARRYB[14][5] ) );
  NAND3X1 U501 ( .A(n891), .B(n890), .C(n892), .Y(n336) );
  XOR2X1 U502 ( .A(n338), .B(n337), .Y(\SUMB[2][9] ) );
  XOR2X1 U503 ( .A(n974), .B(\ab[2][9] ), .Y(n338) );
  XOR2X1 U504 ( .A(\CARRYB[10][3] ), .B(\ab[11][3] ), .Y(n763) );
  XOR2X1 U505 ( .A(n339), .B(n414), .Y(\SUMB[12][4] ) );
  XOR2X1 U506 ( .A(\SUMB[1][3] ), .B(\ab[2][2] ), .Y(n340) );
  XOR2X1 U507 ( .A(n63), .B(n340), .Y(\SUMB[2][2] ) );
  NAND2X1 U508 ( .A(n63), .B(\SUMB[1][3] ), .Y(n341) );
  NAND2X1 U509 ( .A(n63), .B(\ab[2][2] ), .Y(n342) );
  NAND2X1 U510 ( .A(\SUMB[1][3] ), .B(\ab[2][2] ), .Y(n343) );
  NAND3X1 U511 ( .A(n342), .B(n341), .C(n343), .Y(\CARRYB[2][2] ) );
  NAND3X1 U512 ( .A(n851), .B(n850), .C(n852), .Y(n344) );
  BUFX2 U513 ( .A(\CARRYB[13][0] ), .Y(n345) );
  XNOR2X1 U514 ( .A(n346), .B(n347), .Y(\SUMB[5][5] ) );
  XOR2X1 U515 ( .A(\CARRYB[4][5] ), .B(\ab[5][5] ), .Y(n346) );
  INVX2 U516 ( .A(\SUMB[4][6] ), .Y(n347) );
  NAND3X1 U517 ( .A(n875), .B(n876), .C(n877), .Y(n348) );
  NAND3X1 U518 ( .A(n744), .B(n745), .C(n746), .Y(n349) );
  INVX2 U519 ( .A(\SUMB[11][5] ), .Y(n414) );
  XOR2X1 U520 ( .A(\ab[3][14] ), .B(\ab[2][15] ), .Y(n350) );
  XOR2X1 U521 ( .A(n350), .B(\CARRYB[2][14] ), .Y(\SUMB[3][14] ) );
  NAND2X1 U522 ( .A(\CARRYB[2][14] ), .B(\ab[3][14] ), .Y(n351) );
  NAND2X1 U523 ( .A(\CARRYB[2][14] ), .B(\ab[2][15] ), .Y(n352) );
  NAND2X1 U524 ( .A(\ab[3][14] ), .B(\ab[2][15] ), .Y(n353) );
  NAND3X1 U525 ( .A(n352), .B(n351), .C(n353), .Y(\CARRYB[3][14] ) );
  XOR2X1 U526 ( .A(\CARRYB[14][7] ), .B(\ab[15][7] ), .Y(n354) );
  XOR2X1 U527 ( .A(\SUMB[14][8] ), .B(n354), .Y(\SUMB[15][7] ) );
  NAND2X1 U528 ( .A(\SUMB[14][8] ), .B(\CARRYB[14][7] ), .Y(n355) );
  NAND2X1 U529 ( .A(\SUMB[14][8] ), .B(\ab[15][7] ), .Y(n356) );
  NAND2X1 U530 ( .A(\CARRYB[14][7] ), .B(\ab[15][7] ), .Y(n357) );
  NAND3X1 U531 ( .A(n356), .B(n355), .C(n357), .Y(\CARRYB[15][7] ) );
  XOR2X1 U532 ( .A(\CARRYB[11][10] ), .B(\ab[12][10] ), .Y(n358) );
  XOR2X1 U533 ( .A(\SUMB[11][11] ), .B(n358), .Y(\SUMB[12][10] ) );
  NAND2X1 U534 ( .A(\SUMB[11][11] ), .B(\CARRYB[11][10] ), .Y(n359) );
  NAND2X1 U535 ( .A(\SUMB[11][11] ), .B(\ab[12][10] ), .Y(n360) );
  NAND2X1 U536 ( .A(\CARRYB[11][10] ), .B(\ab[12][10] ), .Y(n361) );
  NAND3X1 U537 ( .A(n360), .B(n359), .C(n361), .Y(\CARRYB[12][10] ) );
  XOR2X1 U538 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .Y(n362) );
  XOR2X1 U539 ( .A(n362), .B(\SUMB[7][14] ), .Y(\SUMB[8][13] ) );
  NAND2X1 U540 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .Y(n363) );
  NAND2X1 U541 ( .A(\ab[8][13] ), .B(\SUMB[7][14] ), .Y(n364) );
  NAND2X1 U542 ( .A(\CARRYB[7][13] ), .B(\SUMB[7][14] ), .Y(n365) );
  NAND3X1 U543 ( .A(n363), .B(n364), .C(n365), .Y(\CARRYB[8][13] ) );
  XOR2X1 U544 ( .A(\ab[9][13] ), .B(\SUMB[8][14] ), .Y(n366) );
  XOR2X1 U545 ( .A(n366), .B(\CARRYB[8][13] ), .Y(\SUMB[9][13] ) );
  NAND2X1 U546 ( .A(\ab[9][13] ), .B(\SUMB[8][14] ), .Y(n367) );
  NAND2X1 U547 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .Y(n368) );
  NAND2X1 U548 ( .A(\SUMB[8][14] ), .B(\CARRYB[8][13] ), .Y(n369) );
  NAND3X1 U549 ( .A(n367), .B(n368), .C(n369), .Y(\CARRYB[9][13] ) );
  BUFX2 U550 ( .A(n36), .Y(n370) );
  NAND3X1 U551 ( .A(n753), .B(n754), .C(n752), .Y(n371) );
  XNOR2X1 U552 ( .A(n372), .B(\SUMB[4][4] ), .Y(\SUMB[5][3] ) );
  XOR2X1 U553 ( .A(n949), .B(\ab[5][3] ), .Y(n372) );
  XNOR2X1 U554 ( .A(n931), .B(n373), .Y(\SUMB[8][1] ) );
  XOR2X1 U555 ( .A(n376), .B(n426), .Y(n374) );
  INVX1 U556 ( .A(\SUMB[7][4] ), .Y(n375) );
  XOR2X1 U557 ( .A(n376), .B(n426), .Y(\SUMB[10][4] ) );
  AND2X2 U558 ( .A(n846), .B(B[1]), .Y(\ab[1][1] ) );
  XNOR2X1 U559 ( .A(n449), .B(n377), .Y(\SUMB[10][3] ) );
  INVX2 U560 ( .A(\SUMB[9][4] ), .Y(n377) );
  NAND2X1 U561 ( .A(n528), .B(n78), .Y(n977) );
  NAND3X1 U562 ( .A(n814), .B(n813), .C(n815), .Y(n378) );
  NAND3X1 U563 ( .A(n607), .B(n605), .C(n11), .Y(n379) );
  NAND3X1 U564 ( .A(n781), .B(n782), .C(n783), .Y(n380) );
  NAND3X1 U565 ( .A(n881), .B(n33), .C(n882), .Y(n381) );
  INVX1 U566 ( .A(\CARRYB[2][10] ), .Y(n909) );
  NAND2X1 U567 ( .A(\SUMB[10][5] ), .B(n203), .Y(n382) );
  NAND2X1 U568 ( .A(\SUMB[10][5] ), .B(\ab[11][4] ), .Y(n383) );
  NAND2X1 U569 ( .A(n203), .B(\ab[11][4] ), .Y(n384) );
  NAND3X1 U570 ( .A(n384), .B(n382), .C(n383), .Y(\CARRYB[11][4] ) );
  NAND3X1 U571 ( .A(n899), .B(n900), .C(n901), .Y(n385) );
  NAND3X1 U572 ( .A(n747), .B(n119), .C(n749), .Y(n386) );
  NAND3X1 U573 ( .A(n590), .B(n591), .C(n592), .Y(n387) );
  NAND3X1 U574 ( .A(n784), .B(n785), .C(n786), .Y(n388) );
  INVX1 U575 ( .A(\SUMB[13][3] ), .Y(n425) );
  XOR2X1 U576 ( .A(\CARRYB[10][8] ), .B(\ab[11][8] ), .Y(n389) );
  XOR2X1 U577 ( .A(\SUMB[10][9] ), .B(n389), .Y(\SUMB[11][8] ) );
  NAND2X1 U578 ( .A(\SUMB[10][9] ), .B(\CARRYB[10][8] ), .Y(n390) );
  NAND2X1 U579 ( .A(\SUMB[10][9] ), .B(\ab[11][8] ), .Y(n391) );
  NAND2X1 U580 ( .A(\CARRYB[10][8] ), .B(\ab[11][8] ), .Y(n392) );
  NAND3X1 U581 ( .A(n391), .B(n390), .C(n392), .Y(\CARRYB[11][8] ) );
  NAND3X1 U582 ( .A(n697), .B(n699), .C(n123), .Y(n393) );
  NAND3X1 U583 ( .A(n652), .B(n653), .C(n654), .Y(n394) );
  XNOR2X1 U584 ( .A(n648), .B(n395), .Y(\SUMB[3][4] ) );
  INVX1 U585 ( .A(\SUMB[2][5] ), .Y(n395) );
  BUFX2 U586 ( .A(n1025), .Y(n396) );
  XOR2X1 U587 ( .A(\CARRYB[3][3] ), .B(\ab[4][3] ), .Y(n397) );
  XOR2X1 U588 ( .A(\SUMB[3][4] ), .B(n397), .Y(\SUMB[4][3] ) );
  NAND2X1 U589 ( .A(\SUMB[3][4] ), .B(\CARRYB[3][3] ), .Y(n398) );
  NAND2X1 U590 ( .A(\SUMB[3][4] ), .B(\ab[4][3] ), .Y(n399) );
  NAND2X1 U591 ( .A(\CARRYB[3][3] ), .B(\ab[4][3] ), .Y(n400) );
  NAND3X1 U592 ( .A(n400), .B(n399), .C(n398), .Y(\CARRYB[4][3] ) );
  INVX1 U593 ( .A(\CARRYB[4][3] ), .Y(n949) );
  INVX4 U594 ( .A(A[3]), .Y(n1024) );
  AND2X2 U595 ( .A(n236), .B(B[7]), .Y(n435) );
  XOR2X1 U596 ( .A(\SUMB[3][10] ), .B(n401), .Y(n454) );
  XOR2X1 U597 ( .A(n174), .B(\ab[10][2] ), .Y(n402) );
  XOR2X1 U598 ( .A(\SUMB[9][3] ), .B(n402), .Y(\SUMB[10][2] ) );
  NAND2X1 U599 ( .A(\SUMB[9][3] ), .B(\CARRYB[9][2] ), .Y(n403) );
  NAND2X1 U600 ( .A(\SUMB[9][3] ), .B(\ab[10][2] ), .Y(n404) );
  NAND2X1 U601 ( .A(\CARRYB[9][2] ), .B(\ab[10][2] ), .Y(n405) );
  NAND3X1 U602 ( .A(n404), .B(n403), .C(n405), .Y(\CARRYB[10][2] ) );
  XNOR2X1 U603 ( .A(\ab[1][5] ), .B(n406), .Y(\SUMB[1][5] ) );
  NAND2X1 U604 ( .A(B[6]), .B(n987), .Y(n406) );
  NAND2X1 U605 ( .A(\SUMB[4][12] ), .B(n16), .Y(n407) );
  NAND2X1 U606 ( .A(\SUMB[4][12] ), .B(\ab[5][11] ), .Y(n408) );
  NAND2X1 U607 ( .A(n16), .B(\ab[5][11] ), .Y(n409) );
  NAND3X1 U608 ( .A(n408), .B(n407), .C(n409), .Y(\CARRYB[5][11] ) );
  INVX2 U609 ( .A(\CARRYB[5][6] ), .Y(n445) );
  XOR2X1 U610 ( .A(n410), .B(n534), .Y(\SUMB[8][4] ) );
  INVX1 U611 ( .A(\SUMB[3][9] ), .Y(n411) );
  XNOR2X1 U612 ( .A(\CARRYB[3][8] ), .B(\ab[4][8] ), .Y(n412) );
  NAND3X1 U613 ( .A(n453), .B(n452), .C(n451), .Y(n413) );
  BUFX2 U614 ( .A(n75), .Y(n415) );
  XOR2X1 U615 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .Y(n416) );
  XOR2X1 U616 ( .A(n416), .B(\SUMB[7][13] ), .Y(\SUMB[8][12] ) );
  XOR2X1 U617 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .Y(n417) );
  XOR2X1 U618 ( .A(n417), .B(\SUMB[8][12] ), .Y(\SUMB[9][11] ) );
  NAND2X1 U619 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .Y(n418) );
  NAND2X1 U620 ( .A(\ab[8][12] ), .B(\SUMB[7][13] ), .Y(n419) );
  NAND2X1 U621 ( .A(\CARRYB[7][12] ), .B(\SUMB[7][13] ), .Y(n420) );
  NAND3X1 U622 ( .A(n418), .B(n419), .C(n420), .Y(\CARRYB[8][12] ) );
  NAND2X1 U623 ( .A(\ab[9][11] ), .B(n295), .Y(n421) );
  NAND2X1 U624 ( .A(\ab[9][11] ), .B(\SUMB[8][12] ), .Y(n422) );
  NAND2X1 U625 ( .A(n295), .B(\SUMB[8][12] ), .Y(n423) );
  NAND3X1 U626 ( .A(n421), .B(n422), .C(n423), .Y(\CARRYB[9][11] ) );
  INVX2 U627 ( .A(n986), .Y(n511) );
  XOR2X1 U628 ( .A(\SUMB[12][7] ), .B(n424), .Y(\SUMB[13][6] ) );
  XOR2X1 U629 ( .A(n575), .B(n425), .Y(\SUMB[14][2] ) );
  INVX2 U630 ( .A(\SUMB[9][5] ), .Y(n426) );
  XOR2X1 U631 ( .A(\CARRYB[14][3] ), .B(\ab[15][3] ), .Y(n427) );
  XOR2X1 U632 ( .A(\SUMB[14][4] ), .B(n427), .Y(\SUMB[15][3] ) );
  NAND2X1 U633 ( .A(\SUMB[14][4] ), .B(n275), .Y(n428) );
  NAND2X1 U634 ( .A(\SUMB[14][4] ), .B(\ab[15][3] ), .Y(n429) );
  NAND2X1 U635 ( .A(n275), .B(\ab[15][3] ), .Y(n430) );
  NAND3X1 U636 ( .A(n429), .B(n428), .C(n430), .Y(\CARRYB[15][3] ) );
  INVX1 U637 ( .A(B[7]), .Y(n1004) );
  BUFX2 U638 ( .A(\SUMB[10][1] ), .Y(n432) );
  NAND3X1 U639 ( .A(n630), .B(n629), .C(n631), .Y(n433) );
  XNOR2X1 U640 ( .A(\SUMB[4][3] ), .B(n434), .Y(\SUMB[5][2] ) );
  XNOR2X1 U641 ( .A(\CARRYB[4][2] ), .B(\ab[5][2] ), .Y(n434) );
  NAND2X1 U642 ( .A(\ab[3][8] ), .B(n436), .Y(n437) );
  NAND2X1 U643 ( .A(n218), .B(n126), .Y(n438) );
  NAND2X1 U644 ( .A(n437), .B(n438), .Y(n615) );
  AND2X2 U645 ( .A(B[7]), .B(n511), .Y(n439) );
  BUFX2 U646 ( .A(\SUMB[12][1] ), .Y(n443) );
  NAND2X1 U647 ( .A(n445), .B(\ab[6][6] ), .Y(n446) );
  NAND2X1 U648 ( .A(n444), .B(n193), .Y(n447) );
  NAND2X1 U649 ( .A(n446), .B(n447), .Y(n923) );
  INVX1 U650 ( .A(\ab[6][6] ), .Y(n444) );
  XNOR2X1 U651 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .Y(n448) );
  XOR2X1 U652 ( .A(\SUMB[5][4] ), .B(\ab[6][3] ), .Y(n450) );
  XOR2X1 U653 ( .A(n15), .B(n450), .Y(\SUMB[6][3] ) );
  NAND2X1 U654 ( .A(\SUMB[5][4] ), .B(\CARRYB[5][3] ), .Y(n451) );
  NAND2X1 U655 ( .A(\CARRYB[5][3] ), .B(\ab[6][3] ), .Y(n452) );
  NAND2X1 U656 ( .A(\SUMB[5][4] ), .B(\ab[6][3] ), .Y(n453) );
  NAND3X1 U657 ( .A(n453), .B(n451), .C(n452), .Y(\CARRYB[6][3] ) );
  XNOR2X1 U658 ( .A(n454), .B(n978), .Y(\SUMB[4][9] ) );
  XOR2X1 U659 ( .A(n455), .B(n608), .Y(\SUMB[9][2] ) );
  XNOR2X1 U660 ( .A(\ab[9][2] ), .B(n197), .Y(n455) );
  XOR2X1 U661 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .Y(n456) );
  XOR2X1 U662 ( .A(n456), .B(\SUMB[11][10] ), .Y(\SUMB[12][9] ) );
  XOR2X1 U663 ( .A(n457), .B(\SUMB[12][9] ), .Y(\SUMB[13][8] ) );
  NAND2X1 U664 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .Y(n458) );
  NAND2X1 U665 ( .A(\ab[12][9] ), .B(\SUMB[11][10] ), .Y(n459) );
  NAND2X1 U666 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Y(n460) );
  NAND3X1 U667 ( .A(n458), .B(n459), .C(n460), .Y(\CARRYB[12][9] ) );
  NAND2X1 U668 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .Y(n461) );
  NAND2X1 U669 ( .A(\ab[13][8] ), .B(\SUMB[12][9] ), .Y(n462) );
  NAND2X1 U670 ( .A(\CARRYB[12][8] ), .B(\SUMB[12][9] ), .Y(n463) );
  NAND3X1 U671 ( .A(n461), .B(n462), .C(n463), .Y(\CARRYB[13][8] ) );
  XNOR2X1 U672 ( .A(\ab[0][9] ), .B(n464), .Y(\SUMB[1][8] ) );
  NAND2X1 U673 ( .A(n1007), .B(n514), .Y(n464) );
  NAND2X1 U674 ( .A(\ab[9][9] ), .B(n221), .Y(n465) );
  NAND2X1 U675 ( .A(\SUMB[8][10] ), .B(\ab[9][9] ), .Y(n466) );
  NAND2X1 U676 ( .A(n221), .B(\SUMB[8][10] ), .Y(n467) );
  NAND3X1 U677 ( .A(n465), .B(n466), .C(n467), .Y(\CARRYB[9][9] ) );
  NAND2X1 U678 ( .A(\ab[10][8] ), .B(n349), .Y(n468) );
  NAND2X1 U679 ( .A(\ab[10][8] ), .B(\SUMB[9][9] ), .Y(n469) );
  NAND2X1 U680 ( .A(n349), .B(\SUMB[9][9] ), .Y(n470) );
  NAND3X1 U681 ( .A(n468), .B(n469), .C(n470), .Y(\CARRYB[10][8] ) );
  INVX1 U682 ( .A(n1017), .Y(n1038) );
  XNOR2X1 U683 ( .A(n471), .B(\SUMB[3][13] ), .Y(\SUMB[4][12] ) );
  XOR2X1 U684 ( .A(\ab[4][12] ), .B(n593), .Y(n471) );
  NAND2X1 U685 ( .A(n487), .B(n485), .Y(n472) );
  NAND2X1 U686 ( .A(n243), .B(n473), .Y(n980) );
  INVX4 U687 ( .A(B[13]), .Y(n1016) );
  XNOR2X1 U688 ( .A(n371), .B(\ab[13][1] ), .Y(n474) );
  NAND3X1 U689 ( .A(n12), .B(n88), .C(n637), .Y(n475) );
  BUFX2 U690 ( .A(\CARRYB[4][6] ), .Y(n476) );
  INVX4 U691 ( .A(B[11]), .Y(n1012) );
  XOR2X1 U692 ( .A(\SUMB[4][7] ), .B(\ab[5][6] ), .Y(n477) );
  XOR2X1 U693 ( .A(n477), .B(n476), .Y(\SUMB[5][6] ) );
  NAND2X1 U694 ( .A(\SUMB[4][7] ), .B(\CARRYB[4][6] ), .Y(n478) );
  NAND2X1 U695 ( .A(\CARRYB[4][6] ), .B(\ab[5][6] ), .Y(n479) );
  NAND2X1 U696 ( .A(\ab[5][6] ), .B(\SUMB[4][7] ), .Y(n480) );
  NAND3X1 U697 ( .A(n478), .B(n479), .C(n480), .Y(\CARRYB[5][6] ) );
  NAND2X1 U698 ( .A(\SUMB[14][1] ), .B(n316), .Y(n481) );
  NAND2X1 U699 ( .A(\SUMB[14][1] ), .B(\ab[15][0] ), .Y(n482) );
  NAND2X1 U700 ( .A(n316), .B(\ab[15][0] ), .Y(n483) );
  NAND3X1 U701 ( .A(n483), .B(n481), .C(n482), .Y(\CARRYB[15][0] ) );
  NAND3X1 U702 ( .A(n914), .B(n915), .C(n916), .Y(n484) );
  NAND2X1 U703 ( .A(n93), .B(n53), .Y(n485) );
  NAND2X1 U704 ( .A(n93), .B(\ab[12][3] ), .Y(n486) );
  NAND2X1 U705 ( .A(n53), .B(\ab[12][3] ), .Y(n487) );
  NAND3X1 U706 ( .A(n487), .B(n485), .C(n486), .Y(\CARRYB[12][3] ) );
  NAND3X1 U707 ( .A(n757), .B(n756), .C(n758), .Y(n488) );
  NAND3X1 U708 ( .A(n623), .B(n622), .C(n621), .Y(n489) );
  NAND3X1 U709 ( .A(n948), .B(n947), .C(n946), .Y(n490) );
  NAND3X1 U710 ( .A(n913), .B(n912), .C(n911), .Y(n491) );
  NAND3X1 U711 ( .A(n917), .B(n918), .C(n919), .Y(n492) );
  NAND3X1 U712 ( .A(n579), .B(n580), .C(n581), .Y(n493) );
  NAND3X1 U713 ( .A(n671), .B(n670), .C(n672), .Y(n494) );
  XOR2X1 U714 ( .A(\SUMB[2][2] ), .B(\ab[3][1] ), .Y(n495) );
  XOR2X1 U715 ( .A(\CARRYB[2][1] ), .B(n495), .Y(\SUMB[3][1] ) );
  NAND2X1 U716 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n496) );
  NAND2X1 U717 ( .A(\CARRYB[2][1] ), .B(\ab[3][1] ), .Y(n497) );
  NAND2X1 U718 ( .A(\SUMB[2][2] ), .B(\ab[3][1] ), .Y(n498) );
  NAND3X1 U719 ( .A(n497), .B(n496), .C(n498), .Y(\CARRYB[3][1] ) );
  XOR2X1 U720 ( .A(n370), .B(\ab[14][0] ), .Y(n499) );
  XOR2X1 U721 ( .A(n499), .B(n345), .Y(\A1[12] ) );
  NAND2X1 U722 ( .A(\SUMB[13][1] ), .B(\CARRYB[13][0] ), .Y(n500) );
  NAND2X1 U723 ( .A(\CARRYB[13][0] ), .B(\ab[14][0] ), .Y(n501) );
  NAND2X1 U724 ( .A(\SUMB[13][1] ), .B(\ab[14][0] ), .Y(n502) );
  NAND3X1 U725 ( .A(n501), .B(n500), .C(n502), .Y(\CARRYB[14][0] ) );
  XOR2X1 U726 ( .A(\ab[2][3] ), .B(\SUMB[1][4] ), .Y(n504) );
  XOR2X1 U727 ( .A(n970), .B(n504), .Y(\SUMB[2][3] ) );
  NAND2X1 U728 ( .A(n970), .B(\ab[2][3] ), .Y(n505) );
  NAND2X1 U729 ( .A(n970), .B(\SUMB[1][4] ), .Y(n506) );
  NAND2X1 U730 ( .A(\ab[2][3] ), .B(\SUMB[1][4] ), .Y(n507) );
  NAND3X1 U731 ( .A(n506), .B(n505), .C(n507), .Y(\CARRYB[2][3] ) );
  NAND2X1 U732 ( .A(\SUMB[4][3] ), .B(n145), .Y(n508) );
  NAND2X1 U733 ( .A(\SUMB[4][3] ), .B(\ab[5][2] ), .Y(n509) );
  NAND2X1 U734 ( .A(n145), .B(\ab[5][2] ), .Y(n510) );
  NAND3X1 U735 ( .A(n509), .B(n508), .C(n510), .Y(\CARRYB[5][2] ) );
  INVX1 U736 ( .A(n132), .Y(n1042) );
  XOR2X1 U737 ( .A(n512), .B(n513), .Y(\SUMB[3][7] ) );
  XNOR2X1 U738 ( .A(\ab[3][7] ), .B(n302), .Y(n512) );
  INVX1 U739 ( .A(\SUMB[2][8] ), .Y(n513) );
  XOR2X1 U740 ( .A(\SUMB[3][2] ), .B(\ab[4][1] ), .Y(n515) );
  XOR2X1 U741 ( .A(\CARRYB[3][1] ), .B(n515), .Y(\SUMB[4][1] ) );
  NAND2X1 U742 ( .A(\SUMB[3][2] ), .B(\CARRYB[3][1] ), .Y(n516) );
  NAND2X1 U743 ( .A(\CARRYB[3][1] ), .B(\ab[4][1] ), .Y(n517) );
  NAND2X1 U744 ( .A(\SUMB[3][2] ), .B(\ab[4][1] ), .Y(n518) );
  NAND3X1 U745 ( .A(n517), .B(n516), .C(n518), .Y(\CARRYB[4][1] ) );
  XOR2X1 U746 ( .A(n181), .B(\ab[2][6] ), .Y(n519) );
  NAND2X1 U747 ( .A(\SUMB[1][7] ), .B(n181), .Y(n520) );
  NAND2X1 U748 ( .A(\SUMB[1][7] ), .B(\ab[2][6] ), .Y(n521) );
  NAND2X1 U749 ( .A(n181), .B(\ab[2][6] ), .Y(n522) );
  NAND3X1 U750 ( .A(n520), .B(n521), .C(n522), .Y(\CARRYB[2][6] ) );
  NAND3X1 U751 ( .A(n559), .B(n558), .C(n560), .Y(n523) );
  INVX1 U752 ( .A(n1013), .Y(n1040) );
  AND2X2 U753 ( .A(n999), .B(n514), .Y(n525) );
  BUFX2 U754 ( .A(\SUMB[1][6] ), .Y(n526) );
  INVX1 U755 ( .A(n1009), .Y(n1041) );
  NAND2X1 U756 ( .A(\SUMB[1][10] ), .B(\CARRYB[1][9] ), .Y(n527) );
  NAND2X1 U757 ( .A(\SUMB[1][10] ), .B(\ab[2][9] ), .Y(n528) );
  NAND2X1 U758 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .Y(n529) );
  NAND3X1 U759 ( .A(n528), .B(n527), .C(n529), .Y(\CARRYB[2][9] ) );
  XNOR2X1 U760 ( .A(\CARRYB[13][1] ), .B(n530), .Y(n633) );
  BUFX2 U761 ( .A(\SUMB[6][3] ), .Y(n531) );
  XNOR2X1 U762 ( .A(n532), .B(\SUMB[3][8] ), .Y(\SUMB[4][7] ) );
  NAND3X1 U763 ( .A(n649), .B(n650), .C(n651), .Y(n533) );
  XOR2X1 U764 ( .A(\CARRYB[10][6] ), .B(\ab[11][6] ), .Y(n535) );
  XOR2X1 U765 ( .A(n535), .B(\SUMB[10][7] ), .Y(\SUMB[11][6] ) );
  NAND2X1 U766 ( .A(\SUMB[10][7] ), .B(n379), .Y(n536) );
  NAND2X1 U767 ( .A(\SUMB[10][7] ), .B(\ab[11][6] ), .Y(n537) );
  NAND2X1 U768 ( .A(n379), .B(\ab[11][6] ), .Y(n538) );
  NAND3X1 U769 ( .A(n537), .B(n536), .C(n538), .Y(\CARRYB[11][6] ) );
  NAND3X1 U770 ( .A(n787), .B(n789), .C(n788), .Y(n539) );
  NAND3X1 U771 ( .A(n611), .B(n610), .C(n612), .Y(n540) );
  INVX2 U772 ( .A(n1000), .Y(n985) );
  XNOR2X1 U773 ( .A(n700), .B(n541), .Y(\SUMB[6][5] ) );
  INVX2 U774 ( .A(\SUMB[5][6] ), .Y(n541) );
  INVX1 U775 ( .A(n951), .Y(n939) );
  INVX4 U776 ( .A(B[9]), .Y(n1008) );
  XNOR2X1 U777 ( .A(n543), .B(n247), .Y(\SUMB[5][7] ) );
  NAND2X1 U778 ( .A(\ab[13][7] ), .B(n19), .Y(n544) );
  NAND2X1 U779 ( .A(\SUMB[12][8] ), .B(\ab[13][7] ), .Y(n545) );
  NAND2X1 U780 ( .A(n19), .B(\SUMB[12][8] ), .Y(n546) );
  NAND3X1 U781 ( .A(n544), .B(n545), .C(n546), .Y(\CARRYB[13][7] ) );
  NAND2X1 U782 ( .A(\ab[14][6] ), .B(n393), .Y(n547) );
  NAND2X1 U783 ( .A(\SUMB[13][7] ), .B(\ab[14][6] ), .Y(n548) );
  NAND2X1 U784 ( .A(\SUMB[13][7] ), .B(n393), .Y(n549) );
  NAND3X1 U785 ( .A(n547), .B(n548), .C(n549), .Y(\CARRYB[14][6] ) );
  NAND2X1 U786 ( .A(\SUMB[2][13] ), .B(n238), .Y(n550) );
  NAND2X1 U787 ( .A(\SUMB[2][13] ), .B(\ab[3][12] ), .Y(n551) );
  NAND2X1 U788 ( .A(n238), .B(\ab[3][12] ), .Y(n552) );
  NAND3X1 U789 ( .A(n551), .B(n550), .C(n552), .Y(\CARRYB[3][12] ) );
  XOR2X1 U790 ( .A(\SUMB[9][10] ), .B(\ab[10][9] ), .Y(n553) );
  XOR2X1 U791 ( .A(n553), .B(\CARRYB[9][9] ), .Y(\SUMB[10][9] ) );
  NAND2X1 U792 ( .A(\CARRYB[9][9] ), .B(\SUMB[9][10] ), .Y(n554) );
  NAND2X1 U793 ( .A(\CARRYB[9][9] ), .B(\ab[10][9] ), .Y(n555) );
  NAND2X1 U794 ( .A(\SUMB[9][10] ), .B(\ab[10][9] ), .Y(n556) );
  NAND3X1 U795 ( .A(n555), .B(n554), .C(n556), .Y(\CARRYB[10][9] ) );
  NAND3X1 U796 ( .A(n792), .B(n120), .C(n280), .Y(n557) );
  NAND2X1 U797 ( .A(\CARRYB[3][5] ), .B(\SUMB[3][6] ), .Y(n558) );
  NAND2X1 U798 ( .A(\CARRYB[3][5] ), .B(\ab[4][5] ), .Y(n559) );
  NAND2X1 U799 ( .A(\SUMB[3][6] ), .B(\ab[4][5] ), .Y(n560) );
  NAND3X1 U800 ( .A(n560), .B(n559), .C(n558), .Y(\CARRYB[4][5] ) );
  XOR2X1 U801 ( .A(n561), .B(\SUMB[14][2] ), .Y(\SUMB[15][1] ) );
  NAND2X1 U802 ( .A(\SUMB[14][2] ), .B(n475), .Y(n562) );
  NAND2X1 U803 ( .A(\SUMB[14][2] ), .B(\ab[15][1] ), .Y(n563) );
  NAND2X1 U804 ( .A(n475), .B(\ab[15][1] ), .Y(n564) );
  NAND3X1 U805 ( .A(n564), .B(n562), .C(n563), .Y(\CARRYB[15][1] ) );
  NAND3X1 U806 ( .A(n840), .B(n841), .C(n842), .Y(n565) );
  NAND3X1 U807 ( .A(n634), .B(n636), .C(n635), .Y(n566) );
  NAND2X1 U808 ( .A(\SUMB[5][3] ), .B(\CARRYB[5][2] ), .Y(n567) );
  NAND2X1 U809 ( .A(\CARRYB[5][2] ), .B(\ab[6][2] ), .Y(n568) );
  NAND2X1 U810 ( .A(\SUMB[5][3] ), .B(\ab[6][2] ), .Y(n569) );
  NAND3X1 U811 ( .A(n568), .B(n567), .C(n569), .Y(\CARRYB[6][2] ) );
  XNOR2X1 U812 ( .A(n952), .B(\ab[5][1] ), .Y(n857) );
  INVX1 U813 ( .A(n1015), .Y(n1039) );
  BUFX4 U814 ( .A(\CARRYB[3][9] ), .Y(n978) );
  XNOR2X1 U815 ( .A(n570), .B(\SUMB[12][5] ), .Y(\SUMB[13][4] ) );
  XNOR2X1 U816 ( .A(\CARRYB[12][4] ), .B(\ab[13][4] ), .Y(n570) );
  INVX1 U817 ( .A(n593), .Y(n594) );
  XOR2X1 U818 ( .A(\ab[2][14] ), .B(\ab[1][15] ), .Y(n571) );
  XOR2X1 U819 ( .A(n415), .B(n571), .Y(\SUMB[2][14] ) );
  NAND2X1 U820 ( .A(n75), .B(\ab[2][14] ), .Y(n572) );
  NAND2X1 U821 ( .A(n75), .B(\ab[1][15] ), .Y(n573) );
  NAND2X1 U822 ( .A(\ab[2][14] ), .B(\ab[1][15] ), .Y(n574) );
  NAND3X1 U823 ( .A(n573), .B(n572), .C(n574), .Y(\CARRYB[2][14] ) );
  XNOR2X1 U824 ( .A(n566), .B(\ab[14][2] ), .Y(n575) );
  INVX4 U825 ( .A(B[14]), .Y(n1018) );
  NAND2X1 U826 ( .A(\ab[12][2] ), .B(n492), .Y(n576) );
  NAND2X1 U827 ( .A(n331), .B(\ab[12][2] ), .Y(n577) );
  NAND2X1 U828 ( .A(n331), .B(n492), .Y(n578) );
  NAND3X1 U829 ( .A(n576), .B(n578), .C(n577), .Y(\CARRYB[12][2] ) );
  NAND2X1 U830 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .Y(n579) );
  NAND2X1 U831 ( .A(\SUMB[12][2] ), .B(\ab[13][1] ), .Y(n580) );
  NAND2X1 U832 ( .A(\SUMB[12][2] ), .B(\CARRYB[12][1] ), .Y(n581) );
  NAND3X1 U833 ( .A(n581), .B(n580), .C(n579), .Y(\CARRYB[13][1] ) );
  INVX4 U834 ( .A(n1020), .Y(n987) );
  INVX1 U835 ( .A(n909), .Y(n910) );
  XOR2X1 U836 ( .A(n432), .B(\ab[11][0] ), .Y(n582) );
  XOR2X1 U837 ( .A(n240), .B(n582), .Y(\A1[9] ) );
  NAND2X1 U838 ( .A(\CARRYB[10][0] ), .B(\SUMB[10][1] ), .Y(n583) );
  NAND2X1 U839 ( .A(\CARRYB[10][0] ), .B(\ab[11][0] ), .Y(n584) );
  NAND2X1 U840 ( .A(\SUMB[10][1] ), .B(\ab[11][0] ), .Y(n585) );
  NAND3X1 U841 ( .A(n585), .B(n583), .C(n584), .Y(\CARRYB[11][0] ) );
  NAND2X1 U842 ( .A(\ab[11][7] ), .B(n386), .Y(n587) );
  NAND2X1 U843 ( .A(\SUMB[10][8] ), .B(\ab[11][7] ), .Y(n588) );
  NAND2X1 U844 ( .A(\SUMB[10][8] ), .B(n386), .Y(n589) );
  NAND3X1 U845 ( .A(n587), .B(n588), .C(n589), .Y(\CARRYB[11][7] ) );
  NAND2X1 U846 ( .A(\ab[12][6] ), .B(n279), .Y(n590) );
  NAND2X1 U847 ( .A(\ab[12][6] ), .B(n76), .Y(n591) );
  NAND2X1 U848 ( .A(n279), .B(n76), .Y(n592) );
  NAND3X1 U849 ( .A(n590), .B(n592), .C(n591), .Y(\CARRYB[12][6] ) );
  INVX2 U850 ( .A(\CARRYB[3][12] ), .Y(n593) );
  NAND2X1 U851 ( .A(\SUMB[3][9] ), .B(n565), .Y(n595) );
  NAND2X1 U852 ( .A(\SUMB[3][9] ), .B(\ab[4][8] ), .Y(n596) );
  NAND2X1 U853 ( .A(n565), .B(\ab[4][8] ), .Y(n597) );
  NAND3X1 U854 ( .A(n597), .B(n595), .C(n596), .Y(\CARRYB[4][8] ) );
  XOR2X1 U855 ( .A(\SUMB[10][6] ), .B(n598), .Y(\SUMB[11][5] ) );
  NAND2X1 U856 ( .A(\ab[11][5] ), .B(n276), .Y(n599) );
  NAND2X1 U857 ( .A(\SUMB[10][6] ), .B(\ab[11][5] ), .Y(n600) );
  NAND2X1 U858 ( .A(\SUMB[10][6] ), .B(n276), .Y(n601) );
  NAND3X1 U859 ( .A(n599), .B(n600), .C(n601), .Y(\CARRYB[11][5] ) );
  NAND2X1 U860 ( .A(\ab[12][4] ), .B(n180), .Y(n602) );
  NAND2X1 U861 ( .A(\ab[12][4] ), .B(\SUMB[11][5] ), .Y(n603) );
  NAND2X1 U862 ( .A(\SUMB[11][5] ), .B(n180), .Y(n604) );
  NAND3X1 U863 ( .A(n602), .B(n603), .C(n604), .Y(\CARRYB[12][4] ) );
  NAND2X1 U864 ( .A(\SUMB[9][7] ), .B(n87), .Y(n605) );
  NAND2X1 U865 ( .A(\SUMB[9][7] ), .B(\ab[10][6] ), .Y(n606) );
  NAND2X1 U866 ( .A(n87), .B(\ab[10][6] ), .Y(n607) );
  NAND3X1 U867 ( .A(n607), .B(n605), .C(n606), .Y(\CARRYB[10][6] ) );
  XOR2X1 U868 ( .A(\CARRYB[11][5] ), .B(\ab[12][5] ), .Y(n609) );
  XOR2X1 U869 ( .A(n609), .B(\SUMB[11][6] ), .Y(\SUMB[12][5] ) );
  NAND2X1 U870 ( .A(\SUMB[11][6] ), .B(n328), .Y(n610) );
  NAND2X1 U871 ( .A(\SUMB[11][6] ), .B(\ab[12][5] ), .Y(n611) );
  NAND2X1 U872 ( .A(n328), .B(\ab[12][5] ), .Y(n612) );
  NAND3X1 U873 ( .A(n612), .B(n610), .C(n611), .Y(\CARRYB[12][5] ) );
  NAND3X1 U874 ( .A(n761), .B(n760), .C(n762), .Y(n613) );
  NAND3X1 U875 ( .A(n927), .B(n928), .C(n929), .Y(n614) );
  XOR2X1 U876 ( .A(n443), .B(\ab[13][0] ), .Y(n616) );
  XOR2X1 U877 ( .A(n144), .B(n616), .Y(\A1[11] ) );
  NAND2X1 U878 ( .A(\CARRYB[12][0] ), .B(\SUMB[12][1] ), .Y(n617) );
  NAND2X1 U879 ( .A(\CARRYB[12][0] ), .B(\ab[13][0] ), .Y(n618) );
  NAND2X1 U880 ( .A(\SUMB[12][1] ), .B(\ab[13][0] ), .Y(n619) );
  NAND3X1 U881 ( .A(n619), .B(n617), .C(n618), .Y(\CARRYB[13][0] ) );
  NAND3X1 U882 ( .A(n704), .B(n705), .C(n706), .Y(n620) );
  NAND2X1 U883 ( .A(n980), .B(\ab[13][3] ), .Y(n621) );
  NAND2X1 U884 ( .A(\SUMB[12][4] ), .B(\ab[13][3] ), .Y(n622) );
  NAND2X1 U885 ( .A(n980), .B(\SUMB[12][4] ), .Y(n623) );
  NAND3X1 U886 ( .A(n623), .B(n622), .C(n621), .Y(\CARRYB[13][3] ) );
  NAND2X1 U887 ( .A(\CARRYB[13][2] ), .B(\ab[14][2] ), .Y(n624) );
  NAND2X1 U888 ( .A(\SUMB[13][3] ), .B(\ab[14][2] ), .Y(n625) );
  NAND2X1 U889 ( .A(\CARRYB[13][2] ), .B(\SUMB[13][3] ), .Y(n626) );
  NAND3X1 U890 ( .A(n624), .B(n625), .C(n626), .Y(\CARRYB[14][2] ) );
  NAND2X1 U891 ( .A(n940), .B(n941), .Y(n627) );
  XOR2X1 U892 ( .A(\SUMB[8][2] ), .B(\ab[9][1] ), .Y(n628) );
  XOR2X1 U893 ( .A(n632), .B(n628), .Y(\SUMB[9][1] ) );
  NAND2X1 U894 ( .A(\SUMB[8][2] ), .B(\CARRYB[8][1] ), .Y(n629) );
  NAND2X1 U895 ( .A(\CARRYB[8][1] ), .B(\ab[9][1] ), .Y(n630) );
  NAND2X1 U896 ( .A(\SUMB[8][2] ), .B(\ab[9][1] ), .Y(n631) );
  NAND3X1 U897 ( .A(n631), .B(n629), .C(n630), .Y(\CARRYB[9][1] ) );
  BUFX2 U898 ( .A(\CARRYB[8][1] ), .Y(n632) );
  XOR2X1 U899 ( .A(n633), .B(\SUMB[13][2] ), .Y(\SUMB[14][1] ) );
  NAND2X1 U900 ( .A(\ab[13][2] ), .B(n231), .Y(n634) );
  NAND2X1 U901 ( .A(\ab[13][2] ), .B(\SUMB[12][3] ), .Y(n635) );
  NAND2X1 U902 ( .A(\SUMB[12][3] ), .B(n231), .Y(n636) );
  NAND3X1 U903 ( .A(n634), .B(n636), .C(n635), .Y(\CARRYB[13][2] ) );
  NAND2X1 U904 ( .A(n493), .B(\ab[14][1] ), .Y(n637) );
  NAND2X1 U905 ( .A(\SUMB[13][2] ), .B(\ab[14][1] ), .Y(n638) );
  NAND2X1 U906 ( .A(\SUMB[13][2] ), .B(n493), .Y(n639) );
  NAND3X1 U907 ( .A(n637), .B(n639), .C(n638), .Y(\CARRYB[14][1] ) );
  NOR2X1 U908 ( .A(n1022), .B(n998), .Y(\ab[2][4] ) );
  XOR2X1 U909 ( .A(\ab[4][4] ), .B(n394), .Y(n640) );
  XOR2X1 U910 ( .A(n640), .B(n196), .Y(\SUMB[4][4] ) );
  NAND2X1 U911 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .Y(n641) );
  NAND2X1 U912 ( .A(\ab[4][4] ), .B(\SUMB[3][5] ), .Y(n642) );
  NAND2X1 U913 ( .A(\CARRYB[3][4] ), .B(\SUMB[3][5] ), .Y(n643) );
  NAND2X1 U914 ( .A(\ab[5][3] ), .B(n185), .Y(n644) );
  NAND2X1 U915 ( .A(\SUMB[4][4] ), .B(\ab[5][3] ), .Y(n645) );
  NAND2X1 U916 ( .A(n185), .B(\SUMB[4][4] ), .Y(n646) );
  NAND3X1 U917 ( .A(n645), .B(n644), .C(n646), .Y(\CARRYB[5][3] ) );
  XOR2X1 U918 ( .A(n62), .B(n950), .Y(n647) );
  XOR2X1 U919 ( .A(n647), .B(n526), .Y(\SUMB[2][5] ) );
  XOR2X1 U920 ( .A(\CARRYB[2][4] ), .B(\ab[3][4] ), .Y(n648) );
  NAND2X1 U921 ( .A(n62), .B(n950), .Y(n649) );
  NAND2X1 U922 ( .A(\SUMB[1][6] ), .B(n62), .Y(n650) );
  NAND2X1 U923 ( .A(n950), .B(\SUMB[1][6] ), .Y(n651) );
  NAND3X1 U924 ( .A(n649), .B(n650), .C(n651), .Y(\CARRYB[2][5] ) );
  NAND2X1 U925 ( .A(\CARRYB[2][4] ), .B(\ab[3][4] ), .Y(n652) );
  NAND2X1 U926 ( .A(\ab[3][4] ), .B(\SUMB[2][5] ), .Y(n653) );
  NAND2X1 U927 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n654) );
  NAND3X1 U928 ( .A(n652), .B(n653), .C(n654), .Y(\CARRYB[3][4] ) );
  NAND2X1 U929 ( .A(\SUMB[14][3] ), .B(n202), .Y(n655) );
  NAND2X1 U930 ( .A(\SUMB[14][3] ), .B(\ab[15][2] ), .Y(n656) );
  NAND2X1 U931 ( .A(n202), .B(\ab[15][2] ), .Y(n657) );
  NAND3X1 U932 ( .A(n657), .B(n655), .C(n656), .Y(\CARRYB[15][2] ) );
  NAND2X1 U933 ( .A(\ab[13][4] ), .B(n277), .Y(n658) );
  NAND2X1 U934 ( .A(\SUMB[12][5] ), .B(\ab[13][4] ), .Y(n659) );
  NAND2X1 U935 ( .A(\SUMB[12][5] ), .B(n277), .Y(n660) );
  NAND3X1 U936 ( .A(n658), .B(n659), .C(n660), .Y(\CARRYB[13][4] ) );
  NAND2X1 U937 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .Y(n661) );
  NAND2X1 U938 ( .A(\ab[14][3] ), .B(\SUMB[13][4] ), .Y(n662) );
  NAND2X1 U939 ( .A(\CARRYB[13][3] ), .B(\SUMB[13][4] ), .Y(n663) );
  NAND3X1 U940 ( .A(n663), .B(n661), .C(n662), .Y(\CARRYB[14][3] ) );
  NAND2X1 U941 ( .A(\SUMB[5][5] ), .B(n613), .Y(n664) );
  NAND2X1 U942 ( .A(\SUMB[5][5] ), .B(\ab[6][4] ), .Y(n665) );
  NAND2X1 U943 ( .A(n613), .B(\ab[6][4] ), .Y(n666) );
  NAND2X1 U944 ( .A(n41), .B(n737), .Y(n667) );
  NAND2X1 U945 ( .A(\SUMB[1][9] ), .B(n737), .Y(n668) );
  NAND2X1 U946 ( .A(\SUMB[1][9] ), .B(n41), .Y(n669) );
  NAND3X1 U947 ( .A(n667), .B(n668), .C(n669), .Y(\CARRYB[2][8] ) );
  NAND2X1 U948 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .Y(n670) );
  NAND2X1 U949 ( .A(\SUMB[2][8] ), .B(\ab[3][7] ), .Y(n671) );
  NAND2X1 U950 ( .A(\SUMB[2][8] ), .B(\CARRYB[2][7] ), .Y(n672) );
  NAND3X1 U951 ( .A(n670), .B(n671), .C(n672), .Y(\CARRYB[3][7] ) );
  NAND2X1 U952 ( .A(\SUMB[7][5] ), .B(n620), .Y(n673) );
  NAND2X1 U953 ( .A(\SUMB[7][5] ), .B(\ab[8][4] ), .Y(n674) );
  NAND2X1 U954 ( .A(n620), .B(\ab[8][4] ), .Y(n675) );
  NAND3X1 U955 ( .A(n675), .B(n673), .C(n674), .Y(\CARRYB[8][4] ) );
  XOR2X1 U956 ( .A(\SUMB[14][5] ), .B(n676), .Y(\SUMB[15][4] ) );
  NAND2X1 U957 ( .A(\SUMB[14][5] ), .B(n380), .Y(n677) );
  NAND2X1 U958 ( .A(\SUMB[14][5] ), .B(\ab[15][4] ), .Y(n678) );
  NAND2X1 U959 ( .A(n380), .B(\ab[15][4] ), .Y(n679) );
  XOR2X1 U960 ( .A(n680), .B(\SUMB[6][13] ), .Y(\SUMB[7][12] ) );
  NAND2X1 U961 ( .A(\ab[7][12] ), .B(n713), .Y(n681) );
  NAND2X1 U962 ( .A(\ab[7][12] ), .B(\SUMB[6][13] ), .Y(n682) );
  NAND2X1 U963 ( .A(n713), .B(\SUMB[6][13] ), .Y(n683) );
  NAND3X1 U964 ( .A(n681), .B(n682), .C(n683), .Y(\CARRYB[7][12] ) );
  NAND2X1 U965 ( .A(\ab[8][11] ), .B(n26), .Y(n684) );
  NAND2X1 U966 ( .A(\ab[8][11] ), .B(\SUMB[7][12] ), .Y(n685) );
  NAND2X1 U967 ( .A(n26), .B(\SUMB[7][12] ), .Y(n686) );
  NAND3X1 U968 ( .A(n684), .B(n685), .C(n686), .Y(\CARRYB[8][11] ) );
  XOR2X1 U969 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .Y(n687) );
  XOR2X1 U970 ( .A(n687), .B(\SUMB[4][14] ), .Y(\SUMB[5][13] ) );
  NAND2X1 U971 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .Y(n688) );
  NAND2X1 U972 ( .A(\ab[5][13] ), .B(\SUMB[4][14] ), .Y(n689) );
  NAND2X1 U973 ( .A(\CARRYB[4][13] ), .B(\SUMB[4][14] ), .Y(n690) );
  NAND3X1 U974 ( .A(n688), .B(n689), .C(n690), .Y(\CARRYB[5][13] ) );
  NAND2X1 U975 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .Y(n691) );
  NAND2X1 U976 ( .A(\ab[6][12] ), .B(\SUMB[5][13] ), .Y(n692) );
  NAND2X1 U977 ( .A(\CARRYB[5][12] ), .B(\SUMB[5][13] ), .Y(n693) );
  NAND3X1 U978 ( .A(n691), .B(n692), .C(n693), .Y(\CARRYB[6][12] ) );
  NAND2X1 U979 ( .A(\ab[12][7] ), .B(n124), .Y(n694) );
  NAND2X1 U980 ( .A(\SUMB[11][8] ), .B(\ab[12][7] ), .Y(n695) );
  NAND2X1 U981 ( .A(\SUMB[11][8] ), .B(n124), .Y(n696) );
  NAND3X1 U982 ( .A(n694), .B(n695), .C(n696), .Y(\CARRYB[12][7] ) );
  NAND2X1 U983 ( .A(\ab[13][6] ), .B(n387), .Y(n697) );
  NAND2X1 U984 ( .A(\SUMB[12][7] ), .B(\ab[13][6] ), .Y(n698) );
  NAND2X1 U985 ( .A(\SUMB[12][7] ), .B(n387), .Y(n699) );
  NAND3X1 U986 ( .A(n697), .B(n699), .C(n698), .Y(\CARRYB[13][6] ) );
  NAND2X1 U987 ( .A(n245), .B(\ab[6][5] ), .Y(n701) );
  NAND2X1 U988 ( .A(\ab[6][5] ), .B(\SUMB[5][6] ), .Y(n702) );
  NAND2X1 U989 ( .A(n245), .B(\SUMB[5][6] ), .Y(n703) );
  NAND3X1 U990 ( .A(n701), .B(n702), .C(n703), .Y(\CARRYB[6][5] ) );
  NAND2X1 U991 ( .A(\ab[7][4] ), .B(n122), .Y(n704) );
  NAND2X1 U992 ( .A(\SUMB[6][5] ), .B(\ab[7][4] ), .Y(n705) );
  NAND2X1 U993 ( .A(\SUMB[6][5] ), .B(n122), .Y(n706) );
  NAND3X1 U994 ( .A(n704), .B(n705), .C(n706), .Y(\CARRYB[7][4] ) );
  XOR2X1 U995 ( .A(\CARRYB[2][5] ), .B(\ab[3][5] ), .Y(n707) );
  XOR2X1 U996 ( .A(\SUMB[2][6] ), .B(n707), .Y(\SUMB[3][5] ) );
  NAND2X1 U997 ( .A(\SUMB[2][6] ), .B(n533), .Y(n708) );
  NAND2X1 U998 ( .A(\SUMB[2][6] ), .B(\ab[3][5] ), .Y(n709) );
  NAND2X1 U999 ( .A(n533), .B(\ab[3][5] ), .Y(n710) );
  NAND3X1 U1000 ( .A(n709), .B(n708), .C(n710), .Y(\CARRYB[3][5] ) );
  INVX2 U1001 ( .A(\CARRYB[5][12] ), .Y(n711) );
  INVX2 U1002 ( .A(\CARRYB[6][12] ), .Y(n712) );
  BUFX4 U1003 ( .A(\CARRYB[7][1] ), .Y(n982) );
  NAND2X1 U1004 ( .A(\ab[9][6] ), .B(n442), .Y(n714) );
  NAND2X1 U1005 ( .A(\SUMB[8][7] ), .B(\ab[9][6] ), .Y(n715) );
  NAND2X1 U1006 ( .A(\SUMB[8][7] ), .B(n442), .Y(n716) );
  NAND3X1 U1007 ( .A(n714), .B(n715), .C(n716), .Y(\CARRYB[9][6] ) );
  NAND2X1 U1008 ( .A(n179), .B(\ab[10][5] ), .Y(n717) );
  NAND2X1 U1009 ( .A(\SUMB[9][6] ), .B(n179), .Y(n718) );
  NAND2X1 U1010 ( .A(\SUMB[9][6] ), .B(\ab[10][5] ), .Y(n719) );
  NAND3X1 U1011 ( .A(n717), .B(n718), .C(n719), .Y(\CARRYB[10][5] ) );
  XOR2X1 U1012 ( .A(ZA), .B(ZB), .Y(n720) );
  XOR2X1 U1013 ( .A(n315), .B(n720), .Y(\A1[13] ) );
  NAND2X1 U1014 ( .A(\SUMB[15][0] ), .B(ZA), .Y(n721) );
  NAND2X1 U1015 ( .A(\SUMB[15][0] ), .B(ZB), .Y(n722) );
  NAND2X1 U1016 ( .A(ZA), .B(ZB), .Y(n723) );
  NAND3X1 U1017 ( .A(n723), .B(n721), .C(n722), .Y(\A2[14] ) );
  XNOR2X1 U1018 ( .A(n724), .B(\SUMB[9][2] ), .Y(\SUMB[10][1] ) );
  XNOR2X1 U1019 ( .A(n433), .B(\ab[10][1] ), .Y(n724) );
  XOR2X1 U1020 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .Y(n725) );
  NAND2X1 U1021 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .Y(n727) );
  NAND2X1 U1022 ( .A(\ab[5][10] ), .B(\SUMB[4][11] ), .Y(n728) );
  NAND2X1 U1023 ( .A(\CARRYB[4][10] ), .B(\SUMB[4][11] ), .Y(n729) );
  NAND3X1 U1024 ( .A(n727), .B(n728), .C(n729), .Y(\CARRYB[5][10] ) );
  NAND2X1 U1025 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .Y(n730) );
  NAND2X1 U1026 ( .A(\ab[6][9] ), .B(\SUMB[5][10] ), .Y(n731) );
  NAND2X1 U1027 ( .A(\CARRYB[5][9] ), .B(\SUMB[5][10] ), .Y(n732) );
  NAND3X1 U1028 ( .A(n730), .B(n731), .C(n732), .Y(\CARRYB[6][9] ) );
  NAND2X1 U1029 ( .A(\SUMB[3][12] ), .B(n348), .Y(n733) );
  NAND2X1 U1030 ( .A(\SUMB[3][12] ), .B(\ab[4][11] ), .Y(n734) );
  NAND2X1 U1031 ( .A(n348), .B(\ab[4][11] ), .Y(n735) );
  NAND3X1 U1032 ( .A(n735), .B(n734), .C(n733), .Y(\CARRYB[4][11] ) );
  BUFX2 U1033 ( .A(\CARRYB[4][8] ), .Y(n981) );
  XNOR2X1 U1034 ( .A(n960), .B(\ab[7][2] ), .Y(n930) );
  INVX2 U1035 ( .A(B[1]), .Y(n992) );
  NAND2X1 U1036 ( .A(\ab[3][13] ), .B(n60), .Y(n738) );
  NAND2X1 U1037 ( .A(\ab[3][13] ), .B(\SUMB[2][14] ), .Y(n739) );
  NAND2X1 U1038 ( .A(n60), .B(\SUMB[2][14] ), .Y(n740) );
  NAND3X1 U1039 ( .A(n738), .B(n739), .C(n740), .Y(\CARRYB[3][13] ) );
  NAND2X1 U1040 ( .A(\ab[4][12] ), .B(n594), .Y(n741) );
  NAND2X1 U1041 ( .A(\SUMB[3][13] ), .B(\ab[4][12] ), .Y(n742) );
  NAND2X1 U1042 ( .A(n594), .B(\SUMB[3][13] ), .Y(n743) );
  NAND3X1 U1043 ( .A(n741), .B(n742), .C(n743), .Y(\CARRYB[4][12] ) );
  NAND2X1 U1044 ( .A(\ab[9][8] ), .B(n388), .Y(n744) );
  NAND2X1 U1045 ( .A(\ab[9][8] ), .B(\SUMB[8][9] ), .Y(n745) );
  NAND2X1 U1046 ( .A(n388), .B(\SUMB[8][9] ), .Y(n746) );
  NAND3X1 U1047 ( .A(n744), .B(n745), .C(n746), .Y(\CARRYB[9][8] ) );
  NAND2X1 U1048 ( .A(\ab[10][7] ), .B(n539), .Y(n747) );
  NAND2X1 U1049 ( .A(\ab[10][7] ), .B(\SUMB[9][8] ), .Y(n748) );
  NAND2X1 U1050 ( .A(n539), .B(\SUMB[9][8] ), .Y(n749) );
  NAND3X1 U1051 ( .A(n747), .B(n748), .C(n749), .Y(\CARRYB[10][7] ) );
  XNOR2X1 U1052 ( .A(n750), .B(\SUMB[6][11] ), .Y(\SUMB[7][10] ) );
  XOR2X1 U1053 ( .A(\SUMB[7][3] ), .B(\ab[8][2] ), .Y(n751) );
  XOR2X1 U1054 ( .A(n751), .B(n92), .Y(\SUMB[8][2] ) );
  NAND2X1 U1055 ( .A(\SUMB[11][2] ), .B(\CARRYB[11][1] ), .Y(n752) );
  NAND2X1 U1056 ( .A(\CARRYB[11][1] ), .B(\ab[12][1] ), .Y(n753) );
  NAND2X1 U1057 ( .A(\SUMB[11][2] ), .B(\ab[12][1] ), .Y(n754) );
  NAND3X1 U1058 ( .A(n753), .B(n754), .C(n752), .Y(\CARRYB[12][1] ) );
  NAND2X1 U1059 ( .A(\SUMB[5][8] ), .B(\CARRYB[5][7] ), .Y(n756) );
  NAND2X1 U1060 ( .A(\CARRYB[5][7] ), .B(\ab[6][7] ), .Y(n757) );
  NAND2X1 U1061 ( .A(\SUMB[5][8] ), .B(\ab[6][7] ), .Y(n758) );
  NAND3X1 U1062 ( .A(n758), .B(n756), .C(n757), .Y(\CARRYB[6][7] ) );
  XOR2X1 U1063 ( .A(n260), .B(\ab[5][4] ), .Y(n759) );
  XOR2X1 U1064 ( .A(n121), .B(n759), .Y(\SUMB[5][4] ) );
  NAND2X1 U1065 ( .A(\SUMB[4][5] ), .B(n260), .Y(n760) );
  NAND2X1 U1066 ( .A(\SUMB[4][5] ), .B(\ab[5][4] ), .Y(n761) );
  NAND2X1 U1067 ( .A(n260), .B(\ab[5][4] ), .Y(n762) );
  NAND3X1 U1068 ( .A(n761), .B(n762), .C(n760), .Y(\CARRYB[5][4] ) );
  NAND2X1 U1069 ( .A(\ab[10][4] ), .B(n38), .Y(n764) );
  NAND2X1 U1070 ( .A(\SUMB[9][5] ), .B(\ab[10][4] ), .Y(n765) );
  NAND2X1 U1071 ( .A(\SUMB[9][5] ), .B(n38), .Y(n766) );
  NAND3X1 U1072 ( .A(n764), .B(n765), .C(n766), .Y(\CARRYB[10][4] ) );
  NAND2X1 U1073 ( .A(\ab[11][3] ), .B(n484), .Y(n767) );
  NAND2X1 U1074 ( .A(\ab[11][3] ), .B(\SUMB[10][4] ), .Y(n768) );
  NAND2X1 U1075 ( .A(\SUMB[10][4] ), .B(n484), .Y(n769) );
  NAND3X1 U1076 ( .A(n767), .B(n768), .C(n769), .Y(\CARRYB[11][3] ) );
  XOR2X1 U1077 ( .A(n313), .B(\ab[7][11] ), .Y(n770) );
  XOR2X1 U1078 ( .A(n770), .B(n117), .Y(\SUMB[7][11] ) );
  XOR2X1 U1079 ( .A(\CARRYB[7][10] ), .B(\ab[8][10] ), .Y(n771) );
  XOR2X1 U1080 ( .A(n771), .B(\SUMB[7][11] ), .Y(\SUMB[8][10] ) );
  NAND2X1 U1081 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .Y(n772) );
  NAND2X1 U1082 ( .A(\ab[7][11] ), .B(\SUMB[6][12] ), .Y(n773) );
  NAND2X1 U1083 ( .A(\CARRYB[6][11] ), .B(\SUMB[6][12] ), .Y(n774) );
  NAND3X1 U1084 ( .A(n772), .B(n773), .C(n774), .Y(\CARRYB[7][11] ) );
  NAND2X1 U1085 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .Y(n775) );
  NAND2X1 U1086 ( .A(\ab[8][10] ), .B(\SUMB[7][11] ), .Y(n776) );
  NAND2X1 U1087 ( .A(\CARRYB[7][10] ), .B(\SUMB[7][11] ), .Y(n777) );
  NAND3X1 U1088 ( .A(n775), .B(n776), .C(n777), .Y(\CARRYB[8][10] ) );
  NAND2X1 U1089 ( .A(\ab[13][5] ), .B(n540), .Y(n778) );
  NAND2X1 U1090 ( .A(\SUMB[12][6] ), .B(\ab[13][5] ), .Y(n779) );
  NAND2X1 U1091 ( .A(\SUMB[12][6] ), .B(n540), .Y(n780) );
  NAND3X1 U1092 ( .A(n778), .B(n779), .C(n780), .Y(\CARRYB[13][5] ) );
  NAND2X1 U1093 ( .A(\ab[14][4] ), .B(n330), .Y(n781) );
  NAND2X1 U1094 ( .A(\SUMB[13][5] ), .B(\ab[14][4] ), .Y(n782) );
  NAND2X1 U1095 ( .A(\SUMB[13][5] ), .B(n330), .Y(n783) );
  NAND3X1 U1096 ( .A(n781), .B(n783), .C(n782), .Y(\CARRYB[14][4] ) );
  NAND2X1 U1097 ( .A(\ab[8][8] ), .B(n278), .Y(n784) );
  NAND2X1 U1098 ( .A(\SUMB[7][9] ), .B(\ab[8][8] ), .Y(n785) );
  NAND2X1 U1099 ( .A(n278), .B(\SUMB[7][9] ), .Y(n786) );
  NAND3X1 U1100 ( .A(n784), .B(n785), .C(n786), .Y(\CARRYB[8][8] ) );
  NAND2X1 U1101 ( .A(\ab[9][7] ), .B(n381), .Y(n787) );
  NAND2X1 U1102 ( .A(\SUMB[8][8] ), .B(\ab[9][7] ), .Y(n788) );
  NAND2X1 U1103 ( .A(\SUMB[8][8] ), .B(n381), .Y(n789) );
  NAND3X1 U1104 ( .A(n787), .B(n788), .C(n789), .Y(\CARRYB[9][7] ) );
  XOR2X1 U1105 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .Y(n790) );
  XOR2X1 U1106 ( .A(n790), .B(n95), .Y(\SUMB[6][10] ) );
  XOR2X1 U1107 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .Y(n791) );
  NAND2X1 U1108 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .Y(n792) );
  NAND2X1 U1109 ( .A(\SUMB[5][11] ), .B(\ab[6][10] ), .Y(n793) );
  NAND2X1 U1110 ( .A(\SUMB[5][11] ), .B(\CARRYB[5][10] ), .Y(n794) );
  NAND3X1 U1111 ( .A(n792), .B(n793), .C(n794), .Y(\CARRYB[6][10] ) );
  NAND2X1 U1112 ( .A(\ab[7][9] ), .B(n56), .Y(n795) );
  NAND2X1 U1113 ( .A(\ab[7][9] ), .B(\SUMB[6][10] ), .Y(n796) );
  NAND2X1 U1114 ( .A(n56), .B(\SUMB[6][10] ), .Y(n797) );
  NAND3X1 U1115 ( .A(n795), .B(n796), .C(n797), .Y(\CARRYB[7][9] ) );
  NAND2X1 U1116 ( .A(n811), .B(n79), .Y(n979) );
  NAND2X1 U1117 ( .A(\SUMB[10][2] ), .B(n84), .Y(n798) );
  NAND2X1 U1118 ( .A(\SUMB[10][2] ), .B(\ab[11][1] ), .Y(n799) );
  NAND2X1 U1119 ( .A(n84), .B(\ab[11][1] ), .Y(n800) );
  NAND3X1 U1120 ( .A(n799), .B(n800), .C(n798), .Y(\CARRYB[11][1] ) );
  NAND2X1 U1121 ( .A(\SUMB[6][4] ), .B(\CARRYB[6][3] ), .Y(n801) );
  NAND2X1 U1122 ( .A(\SUMB[6][4] ), .B(\ab[7][3] ), .Y(n802) );
  NAND2X1 U1123 ( .A(\CARRYB[6][3] ), .B(\ab[7][3] ), .Y(n803) );
  NAND3X1 U1124 ( .A(n803), .B(n802), .C(n801), .Y(\CARRYB[7][3] ) );
  NAND2X1 U1125 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .Y(n804) );
  NAND2X1 U1126 ( .A(\ab[6][11] ), .B(\SUMB[5][12] ), .Y(n805) );
  NAND2X1 U1127 ( .A(\CARRYB[5][11] ), .B(\SUMB[5][12] ), .Y(n806) );
  NAND3X1 U1128 ( .A(n804), .B(n805), .C(n806), .Y(\CARRYB[6][11] ) );
  NAND2X1 U1129 ( .A(\ab[7][10] ), .B(n557), .Y(n807) );
  NAND2X1 U1130 ( .A(\ab[7][10] ), .B(\SUMB[6][11] ), .Y(n808) );
  NAND2X1 U1131 ( .A(\SUMB[6][11] ), .B(n557), .Y(n809) );
  NAND3X1 U1132 ( .A(n807), .B(n808), .C(n809), .Y(\CARRYB[7][10] ) );
  NAND2X1 U1133 ( .A(n173), .B(\SUMB[7][4] ), .Y(n810) );
  NAND2X1 U1134 ( .A(\SUMB[7][4] ), .B(\ab[8][3] ), .Y(n811) );
  NAND2X1 U1135 ( .A(n173), .B(\ab[8][3] ), .Y(n812) );
  NAND3X1 U1136 ( .A(n811), .B(n812), .C(n810), .Y(\CARRYB[8][3] ) );
  INVX2 U1137 ( .A(A[1]), .Y(n986) );
  NAND2X1 U1138 ( .A(\SUMB[3][10] ), .B(n978), .Y(n813) );
  NAND2X1 U1139 ( .A(n978), .B(\ab[4][9] ), .Y(n814) );
  NAND2X1 U1140 ( .A(\SUMB[3][10] ), .B(\ab[4][9] ), .Y(n815) );
  NAND3X1 U1141 ( .A(n814), .B(n813), .C(n815), .Y(\CARRYB[4][9] ) );
  NAND2X1 U1142 ( .A(\SUMB[1][11] ), .B(n77), .Y(n816) );
  NAND2X1 U1143 ( .A(n77), .B(\ab[2][10] ), .Y(n817) );
  NAND2X1 U1144 ( .A(\SUMB[1][11] ), .B(\ab[2][10] ), .Y(n818) );
  NAND3X1 U1145 ( .A(n817), .B(n816), .C(n818), .Y(\CARRYB[2][10] ) );
  NAND2X1 U1146 ( .A(\ab[4][6] ), .B(n246), .Y(n819) );
  NAND2X1 U1147 ( .A(\SUMB[3][7] ), .B(\ab[4][6] ), .Y(n820) );
  NAND2X1 U1148 ( .A(n246), .B(\SUMB[3][7] ), .Y(n821) );
  NAND3X1 U1149 ( .A(n819), .B(n820), .C(n821), .Y(\CARRYB[4][6] ) );
  NAND2X1 U1150 ( .A(\ab[5][5] ), .B(n523), .Y(n822) );
  NAND2X1 U1151 ( .A(\SUMB[4][6] ), .B(\ab[5][5] ), .Y(n823) );
  NAND2X1 U1152 ( .A(\SUMB[4][6] ), .B(n523), .Y(n824) );
  NAND3X1 U1153 ( .A(n824), .B(n822), .C(n823), .Y(\CARRYB[5][5] ) );
  NAND2X1 U1154 ( .A(n435), .B(n61), .Y(n825) );
  NAND2X1 U1155 ( .A(\SUMB[1][8] ), .B(n435), .Y(n826) );
  NAND2X1 U1156 ( .A(n61), .B(\SUMB[1][8] ), .Y(n827) );
  NAND3X1 U1157 ( .A(n825), .B(n826), .C(n827), .Y(\CARRYB[2][7] ) );
  NAND2X1 U1158 ( .A(n848), .B(\ab[3][6] ), .Y(n828) );
  NAND2X1 U1159 ( .A(\SUMB[2][7] ), .B(\ab[3][6] ), .Y(n829) );
  NAND2X1 U1160 ( .A(n848), .B(\SUMB[2][7] ), .Y(n830) );
  NAND3X1 U1161 ( .A(n829), .B(n828), .C(n830), .Y(\CARRYB[3][6] ) );
  NAND2X1 U1162 ( .A(\SUMB[6][6] ), .B(\CARRYB[6][5] ), .Y(n831) );
  NAND2X1 U1163 ( .A(\CARRYB[6][5] ), .B(\ab[7][5] ), .Y(n832) );
  NAND2X1 U1164 ( .A(\SUMB[6][6] ), .B(\ab[7][5] ), .Y(n833) );
  NAND3X1 U1165 ( .A(n832), .B(n831), .C(n833), .Y(\CARRYB[7][5] ) );
  NAND2X1 U1166 ( .A(\ab[8][5] ), .B(n303), .Y(n834) );
  NAND2X1 U1167 ( .A(\SUMB[7][6] ), .B(\ab[8][5] ), .Y(n835) );
  NAND2X1 U1168 ( .A(\SUMB[7][6] ), .B(n303), .Y(n836) );
  NAND3X1 U1169 ( .A(n834), .B(n835), .C(n836), .Y(\CARRYB[8][5] ) );
  NAND2X1 U1170 ( .A(n98), .B(\ab[9][4] ), .Y(n837) );
  NAND2X1 U1171 ( .A(\SUMB[8][5] ), .B(n98), .Y(n838) );
  NAND2X1 U1172 ( .A(\SUMB[8][5] ), .B(\ab[9][4] ), .Y(n839) );
  NAND3X1 U1173 ( .A(n837), .B(n839), .C(n838), .Y(\CARRYB[9][4] ) );
  NAND2X1 U1174 ( .A(\ab[3][8] ), .B(n126), .Y(n840) );
  NAND2X1 U1175 ( .A(\SUMB[2][9] ), .B(\ab[3][8] ), .Y(n841) );
  NAND2X1 U1176 ( .A(\SUMB[2][9] ), .B(n126), .Y(n842) );
  NAND3X1 U1177 ( .A(n840), .B(n841), .C(n842), .Y(\CARRYB[3][8] ) );
  NAND2X1 U1178 ( .A(\ab[4][7] ), .B(n494), .Y(n843) );
  NAND2X1 U1179 ( .A(\SUMB[3][8] ), .B(\ab[4][7] ), .Y(n844) );
  NAND2X1 U1180 ( .A(\SUMB[3][8] ), .B(n494), .Y(n845) );
  NAND3X1 U1181 ( .A(n843), .B(n844), .C(n845), .Y(\CARRYB[4][7] ) );
  INVX2 U1182 ( .A(\CARRYB[2][6] ), .Y(n847) );
  XOR2X1 U1183 ( .A(n164), .B(\ab[9][0] ), .Y(n849) );
  XOR2X1 U1184 ( .A(\CARRYB[8][0] ), .B(n849), .Y(\A1[7] ) );
  NAND2X1 U1185 ( .A(\SUMB[8][1] ), .B(\CARRYB[8][0] ), .Y(n850) );
  NAND2X1 U1186 ( .A(\CARRYB[8][0] ), .B(\ab[9][0] ), .Y(n851) );
  NAND2X1 U1187 ( .A(\SUMB[8][1] ), .B(\ab[9][0] ), .Y(n852) );
  NAND3X1 U1188 ( .A(n851), .B(n850), .C(n852), .Y(\CARRYB[9][0] ) );
  XOR2X1 U1189 ( .A(n344), .B(\ab[10][0] ), .Y(n853) );
  XOR2X1 U1190 ( .A(n89), .B(n853), .Y(\A1[8] ) );
  NAND2X1 U1191 ( .A(\SUMB[9][1] ), .B(\CARRYB[9][0] ), .Y(n854) );
  NAND2X1 U1192 ( .A(\SUMB[9][1] ), .B(\ab[10][0] ), .Y(n855) );
  NAND2X1 U1193 ( .A(\CARRYB[9][0] ), .B(\ab[10][0] ), .Y(n856) );
  NAND3X1 U1194 ( .A(n855), .B(n856), .C(n854), .Y(\CARRYB[10][0] ) );
  XOR2X1 U1195 ( .A(n857), .B(\SUMB[4][2] ), .Y(\SUMB[5][1] ) );
  NAND2X1 U1196 ( .A(\SUMB[4][2] ), .B(\CARRYB[4][1] ), .Y(n858) );
  NAND2X1 U1197 ( .A(\SUMB[4][2] ), .B(\ab[5][1] ), .Y(n859) );
  NAND2X1 U1198 ( .A(\CARRYB[4][1] ), .B(\ab[5][1] ), .Y(n860) );
  NAND3X1 U1199 ( .A(n859), .B(n858), .C(n860), .Y(\CARRYB[5][1] ) );
  XOR2X1 U1200 ( .A(\ab[7][0] ), .B(n989), .Y(n861) );
  XOR2X1 U1201 ( .A(n861), .B(\SUMB[6][1] ), .Y(\A1[5] ) );
  NAND2X1 U1202 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .Y(n862) );
  NAND2X1 U1203 ( .A(\ab[6][1] ), .B(\SUMB[5][2] ), .Y(n863) );
  NAND2X1 U1204 ( .A(\CARRYB[5][1] ), .B(\SUMB[5][2] ), .Y(n864) );
  NAND3X1 U1205 ( .A(n862), .B(n863), .C(n864), .Y(\CARRYB[6][1] ) );
  NAND2X1 U1206 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .Y(n865) );
  NAND2X1 U1207 ( .A(\ab[7][0] ), .B(\SUMB[6][1] ), .Y(n866) );
  NAND2X1 U1208 ( .A(\CARRYB[6][0] ), .B(\SUMB[6][1] ), .Y(n867) );
  NAND3X1 U1209 ( .A(n865), .B(n866), .C(n867), .Y(\CARRYB[7][0] ) );
  XOR2X1 U1210 ( .A(\CARRYB[3][2] ), .B(\ab[4][2] ), .Y(n868) );
  XOR2X1 U1211 ( .A(n627), .B(n868), .Y(\SUMB[4][2] ) );
  NAND2X1 U1212 ( .A(\SUMB[3][3] ), .B(n190), .Y(n869) );
  NAND2X1 U1213 ( .A(\SUMB[3][3] ), .B(\ab[4][2] ), .Y(n870) );
  NAND2X1 U1214 ( .A(n190), .B(\ab[4][2] ), .Y(n871) );
  NAND3X1 U1215 ( .A(n870), .B(n869), .C(n871), .Y(\CARRYB[4][2] ) );
  NAND2X1 U1216 ( .A(\CARRYB[1][12] ), .B(\ab[2][12] ), .Y(n872) );
  NAND2X1 U1217 ( .A(\CARRYB[1][12] ), .B(\SUMB[1][13] ), .Y(n873) );
  NAND2X1 U1218 ( .A(\ab[2][12] ), .B(\SUMB[1][13] ), .Y(n874) );
  NAND3X1 U1219 ( .A(n872), .B(n873), .C(n874), .Y(\CARRYB[2][12] ) );
  NAND2X1 U1220 ( .A(\ab[3][11] ), .B(n385), .Y(n875) );
  NAND2X1 U1221 ( .A(\SUMB[2][12] ), .B(\ab[3][11] ), .Y(n876) );
  NAND2X1 U1222 ( .A(\SUMB[2][12] ), .B(n385), .Y(n877) );
  NAND3X1 U1223 ( .A(n875), .B(n876), .C(n877), .Y(\CARRYB[3][11] ) );
  NAND2X1 U1224 ( .A(\ab[7][8] ), .B(n299), .Y(n878) );
  NAND2X1 U1225 ( .A(\SUMB[6][9] ), .B(\ab[7][8] ), .Y(n879) );
  NAND2X1 U1226 ( .A(\SUMB[6][9] ), .B(n299), .Y(n880) );
  NAND3X1 U1227 ( .A(n878), .B(n879), .C(n880), .Y(\CARRYB[7][8] ) );
  NAND2X1 U1228 ( .A(\ab[8][7] ), .B(n329), .Y(n881) );
  NAND2X1 U1229 ( .A(\SUMB[7][8] ), .B(\ab[8][7] ), .Y(n882) );
  NAND2X1 U1230 ( .A(\SUMB[7][8] ), .B(n329), .Y(n883) );
  NAND3X1 U1231 ( .A(n881), .B(n882), .C(n883), .Y(\CARRYB[8][7] ) );
  NAND2X1 U1232 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .Y(n884) );
  NAND2X1 U1233 ( .A(\SUMB[8][3] ), .B(\ab[9][2] ), .Y(n885) );
  NAND2X1 U1234 ( .A(\CARRYB[8][2] ), .B(\SUMB[8][3] ), .Y(n886) );
  NAND3X1 U1235 ( .A(n885), .B(n884), .C(n886), .Y(\CARRYB[9][2] ) );
  NAND2X1 U1236 ( .A(\CARRYB[9][1] ), .B(\ab[10][1] ), .Y(n887) );
  NAND2X1 U1237 ( .A(\SUMB[9][2] ), .B(\CARRYB[9][1] ), .Y(n888) );
  NAND2X1 U1238 ( .A(\ab[10][1] ), .B(\SUMB[9][2] ), .Y(n889) );
  NAND3X1 U1239 ( .A(n887), .B(n888), .C(n889), .Y(\CARRYB[10][1] ) );
  NAND2X1 U1240 ( .A(\SUMB[4][10] ), .B(n378), .Y(n890) );
  NAND2X1 U1241 ( .A(\SUMB[4][10] ), .B(\ab[5][9] ), .Y(n891) );
  NAND2X1 U1242 ( .A(n378), .B(\ab[5][9] ), .Y(n892) );
  NAND3X1 U1243 ( .A(n891), .B(n892), .C(n890), .Y(\CARRYB[5][9] ) );
  NAND2X1 U1244 ( .A(\ab[6][8] ), .B(n490), .Y(n893) );
  NAND2X1 U1245 ( .A(\SUMB[5][9] ), .B(\ab[6][8] ), .Y(n894) );
  NAND2X1 U1246 ( .A(\SUMB[5][9] ), .B(n490), .Y(n895) );
  NAND3X1 U1247 ( .A(n893), .B(n894), .C(n895), .Y(\CARRYB[6][8] ) );
  NAND2X1 U1248 ( .A(\ab[7][7] ), .B(n488), .Y(n896) );
  NAND2X1 U1249 ( .A(\SUMB[6][8] ), .B(\ab[7][7] ), .Y(n897) );
  NAND2X1 U1250 ( .A(\SUMB[6][8] ), .B(n488), .Y(n898) );
  NAND3X1 U1251 ( .A(n896), .B(n897), .C(n898), .Y(\CARRYB[7][7] ) );
  NAND2X1 U1252 ( .A(n222), .B(\ab[2][11] ), .Y(n899) );
  NAND2X1 U1253 ( .A(n222), .B(\SUMB[1][12] ), .Y(n900) );
  NAND2X1 U1254 ( .A(\ab[2][11] ), .B(\SUMB[1][12] ), .Y(n901) );
  NAND3X1 U1255 ( .A(n899), .B(n900), .C(n901), .Y(\CARRYB[2][11] ) );
  NAND2X1 U1256 ( .A(\ab[3][10] ), .B(n910), .Y(n902) );
  NAND2X1 U1257 ( .A(n223), .B(\ab[3][10] ), .Y(n903) );
  NAND2X1 U1258 ( .A(n223), .B(n910), .Y(n904) );
  NAND3X1 U1259 ( .A(n902), .B(n904), .C(n903), .Y(\CARRYB[3][10] ) );
  INVX2 U1260 ( .A(\CARRYB[3][0] ), .Y(n905) );
  INVX4 U1261 ( .A(n905), .Y(n906) );
  INVX2 U1262 ( .A(\CARRYB[4][0] ), .Y(n907) );
  INVX4 U1263 ( .A(n907), .Y(n908) );
  NAND2X1 U1264 ( .A(\SUMB[8][4] ), .B(n979), .Y(n911) );
  NAND2X1 U1265 ( .A(\SUMB[8][4] ), .B(\ab[9][3] ), .Y(n912) );
  NAND2X1 U1266 ( .A(n979), .B(\ab[9][3] ), .Y(n913) );
  NAND3X1 U1267 ( .A(n913), .B(n912), .C(n911), .Y(\CARRYB[9][3] ) );
  NAND2X1 U1268 ( .A(n491), .B(\ab[10][3] ), .Y(n914) );
  NAND2X1 U1269 ( .A(\SUMB[9][4] ), .B(\ab[10][3] ), .Y(n915) );
  NAND2X1 U1270 ( .A(\SUMB[9][4] ), .B(n491), .Y(n916) );
  NAND3X1 U1271 ( .A(n914), .B(n915), .C(n916), .Y(\CARRYB[10][3] ) );
  NAND2X1 U1272 ( .A(n85), .B(\ab[11][2] ), .Y(n917) );
  NAND2X1 U1273 ( .A(\SUMB[10][3] ), .B(\ab[11][2] ), .Y(n918) );
  NAND2X1 U1274 ( .A(\SUMB[10][3] ), .B(n85), .Y(n919) );
  NAND3X1 U1275 ( .A(n917), .B(n918), .C(n919), .Y(\CARRYB[11][2] ) );
  NAND2X1 U1276 ( .A(\SUMB[2][10] ), .B(n977), .Y(n920) );
  NAND2X1 U1277 ( .A(\SUMB[2][10] ), .B(\ab[3][9] ), .Y(n921) );
  NAND2X1 U1278 ( .A(n977), .B(\ab[3][9] ), .Y(n922) );
  NAND3X1 U1279 ( .A(n922), .B(n920), .C(n921), .Y(\CARRYB[3][9] ) );
  XOR2X1 U1280 ( .A(n923), .B(\SUMB[5][7] ), .Y(\SUMB[6][6] ) );
  NAND2X1 U1281 ( .A(\ab[5][7] ), .B(n270), .Y(n924) );
  NAND2X1 U1282 ( .A(n247), .B(\ab[5][7] ), .Y(n925) );
  NAND2X1 U1283 ( .A(n247), .B(n270), .Y(n926) );
  NAND3X1 U1284 ( .A(n924), .B(n925), .C(n926), .Y(\CARRYB[5][7] ) );
  NAND2X1 U1285 ( .A(n193), .B(\ab[6][6] ), .Y(n927) );
  NAND2X1 U1286 ( .A(\SUMB[5][7] ), .B(\ab[6][6] ), .Y(n928) );
  NAND2X1 U1287 ( .A(\SUMB[5][7] ), .B(n230), .Y(n929) );
  NAND3X1 U1288 ( .A(n927), .B(n929), .C(n928), .Y(\CARRYB[6][6] ) );
  XOR2X1 U1289 ( .A(n930), .B(n531), .Y(\SUMB[7][2] ) );
  XOR2X1 U1290 ( .A(\ab[8][1] ), .B(n982), .Y(n931) );
  NAND2X1 U1291 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .Y(n932) );
  NAND2X1 U1292 ( .A(\ab[7][2] ), .B(\SUMB[6][3] ), .Y(n933) );
  NAND2X1 U1293 ( .A(\CARRYB[6][2] ), .B(\SUMB[6][3] ), .Y(n934) );
  NAND3X1 U1294 ( .A(n932), .B(n933), .C(n934), .Y(\CARRYB[7][2] ) );
  NAND2X1 U1295 ( .A(\ab[8][1] ), .B(n982), .Y(n935) );
  NAND2X1 U1296 ( .A(\ab[8][1] ), .B(\SUMB[7][2] ), .Y(n936) );
  NAND2X1 U1297 ( .A(n982), .B(\SUMB[7][2] ), .Y(n937) );
  NAND3X1 U1298 ( .A(n936), .B(n935), .C(n937), .Y(\CARRYB[8][1] ) );
  NAND2X1 U1299 ( .A(\CARRYB[2][3] ), .B(n951), .Y(n940) );
  NAND2X1 U1300 ( .A(n938), .B(n939), .Y(n941) );
  NAND2X1 U1301 ( .A(n940), .B(n941), .Y(\SUMB[3][3] ) );
  INVX1 U1302 ( .A(\CARRYB[2][3] ), .Y(n938) );
  NAND2X1 U1303 ( .A(\SUMB[6][7] ), .B(n614), .Y(n942) );
  NAND2X1 U1304 ( .A(\SUMB[6][7] ), .B(\ab[7][6] ), .Y(n943) );
  NAND2X1 U1305 ( .A(n614), .B(\ab[7][6] ), .Y(n944) );
  NAND3X1 U1306 ( .A(n944), .B(n943), .C(n942), .Y(\CARRYB[7][6] ) );
  XOR2X1 U1307 ( .A(\CARRYB[4][8] ), .B(\ab[5][8] ), .Y(n945) );
  XOR2X1 U1308 ( .A(\SUMB[4][9] ), .B(n945), .Y(\SUMB[5][8] ) );
  NAND2X1 U1309 ( .A(\SUMB[4][9] ), .B(n981), .Y(n946) );
  NAND2X1 U1310 ( .A(\SUMB[4][9] ), .B(\ab[5][8] ), .Y(n947) );
  NAND2X1 U1311 ( .A(n981), .B(\ab[5][8] ), .Y(n948) );
  NAND3X1 U1312 ( .A(n948), .B(n947), .C(n946), .Y(\CARRYB[5][8] ) );
  AND2X2 U1313 ( .A(n524), .B(\ab[1][5] ), .Y(n950) );
  INVX4 U1314 ( .A(A[2]), .Y(n1022) );
  XNOR2X1 U1315 ( .A(\SUMB[2][4] ), .B(\ab[3][3] ), .Y(n951) );
  INVX2 U1316 ( .A(\CARRYB[4][1] ), .Y(n952) );
  XOR2X1 U1317 ( .A(\CARRYB[2][2] ), .B(\ab[3][2] ), .Y(n953) );
  XOR2X1 U1318 ( .A(\SUMB[2][3] ), .B(n953), .Y(\SUMB[3][2] ) );
  NAND2X1 U1319 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(n954) );
  NAND2X1 U1320 ( .A(\SUMB[2][3] ), .B(\ab[3][2] ), .Y(n955) );
  NAND2X1 U1321 ( .A(\CARRYB[2][2] ), .B(\ab[3][2] ), .Y(n956) );
  NAND3X1 U1322 ( .A(n955), .B(n954), .C(n956), .Y(\CARRYB[3][2] ) );
  NAND2X1 U1323 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(n957) );
  NAND2X1 U1324 ( .A(\CARRYB[7][2] ), .B(\ab[8][2] ), .Y(n958) );
  NAND2X1 U1325 ( .A(\SUMB[7][3] ), .B(\ab[8][2] ), .Y(n959) );
  NAND3X1 U1326 ( .A(n959), .B(n957), .C(n958), .Y(\CARRYB[8][2] ) );
  NAND2X1 U1327 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n961) );
  NAND2X1 U1328 ( .A(\CARRYB[2][3] ), .B(\ab[3][3] ), .Y(n962) );
  NAND2X1 U1329 ( .A(\ab[3][3] ), .B(\SUMB[2][4] ), .Y(n963) );
  NAND3X1 U1330 ( .A(n962), .B(n963), .C(n961), .Y(\CARRYB[3][3] ) );
  AND2X2 U1331 ( .A(\CARRYB[15][0] ), .B(\SUMB[15][1] ), .Y(n972) );
  AND2X2 U1332 ( .A(n1025), .B(n1009), .Y(\ab[3][9] ) );
  NOR2X1 U1333 ( .A(n1021), .B(n994), .Y(n964) );
  INVX1 U1334 ( .A(\CARRYB[6][0] ), .Y(n988) );
  AND2X2 U1335 ( .A(\ab[0][5] ), .B(n525), .Y(n965) );
  AND2X2 U1336 ( .A(n228), .B(\CARRYB[15][4] ), .Y(n968) );
  AND2X2 U1337 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n969) );
  AND2X2 U1338 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(n970) );
  AND2X2 U1339 ( .A(\SUMB[15][6] ), .B(\CARRYB[15][5] ), .Y(n973) );
  INVX4 U1340 ( .A(n992), .Y(n993) );
  INVX2 U1341 ( .A(n988), .Y(n989) );
  INVX2 U1342 ( .A(B[0]), .Y(n990) );
  INVX2 U1343 ( .A(A[13]), .Y(n1052) );
  INVX2 U1344 ( .A(ZA), .Y(n1050) );
  INVX2 U1345 ( .A(A[14]), .Y(n1051) );
  INVX2 U1346 ( .A(A[4]), .Y(n1026) );
  INVX2 U1347 ( .A(A[6]), .Y(n1030) );
  INVX2 U1348 ( .A(A[5]), .Y(n1028) );
  INVX2 U1349 ( .A(A[8]), .Y(n1034) );
  INVX2 U1350 ( .A(A[7]), .Y(n1032) );
  INVX2 U1351 ( .A(A[9]), .Y(n1036) );
  XOR2X1 U1352 ( .A(\CARRYB[15][0] ), .B(\SUMB[15][1] ), .Y(\A1[14] ) );
  XOR2X1 U1353 ( .A(\CARRYB[15][1] ), .B(\SUMB[15][2] ), .Y(\A1[15] ) );
  XOR2X1 U1354 ( .A(\SUMB[15][3] ), .B(\CARRYB[15][2] ), .Y(\A1[16] ) );
  XOR2X1 U1355 ( .A(\SUMB[15][4] ), .B(\CARRYB[15][3] ), .Y(\A1[17] ) );
  XOR2X1 U1356 ( .A(\SUMB[15][7] ), .B(\CARRYB[15][6] ), .Y(\A1[20] ) );
  XOR2X1 U1357 ( .A(\SUMB[15][8] ), .B(\CARRYB[15][7] ), .Y(\A1[21] ) );
  XOR2X1 U1358 ( .A(\SUMB[15][9] ), .B(\CARRYB[15][8] ), .Y(\A1[22] ) );
  XOR2X1 U1359 ( .A(\SUMB[15][10] ), .B(\CARRYB[15][9] ), .Y(\A1[23] ) );
  XOR2X1 U1360 ( .A(\SUMB[15][11] ), .B(\CARRYB[15][10] ), .Y(\A1[24] ) );
  XOR2X1 U1361 ( .A(\SUMB[15][12] ), .B(\CARRYB[15][11] ), .Y(\A1[25] ) );
  XOR2X1 U1362 ( .A(\SUMB[15][13] ), .B(\CARRYB[15][12] ), .Y(\A1[26] ) );
  XOR2X1 U1363 ( .A(\SUMB[15][14] ), .B(\CARRYB[15][13] ), .Y(\A1[27] ) );
  XOR2X1 U1364 ( .A(\SUMB[15][15] ), .B(\CARRYB[15][14] ), .Y(\A1[28] ) );
  XOR2X1 U1365 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U1366 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U1367 ( .A(n964), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U1368 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U1369 ( .A(\ab[0][5] ), .B(n525), .Y(\SUMB[1][4] ) );
  XOR2X1 U1370 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U1371 ( .A(n439), .B(\ab[0][8] ), .Y(\SUMB[1][7] ) );
  NAND2X1 U1372 ( .A(n184), .B(\ab[0][10] ), .Y(n974) );
  XOR2X1 U1373 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(\SUMB[1][10] ) );
  XOR2X1 U1374 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Y(\SUMB[1][12] ) );
  NAND2X1 U1375 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Y(n975) );
  XOR2X1 U1376 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Y(\SUMB[1][13] ) );
  NAND2X1 U1377 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Y(n976) );
  INVX2 U1378 ( .A(n976), .Y(\CARRYB[1][13] ) );
  XOR2X1 U1379 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Y(\SUMB[1][14] ) );
  INVX2 U1380 ( .A(n996), .Y(n997) );
  INVX2 U1381 ( .A(n998), .Y(n999) );
  INVX2 U1382 ( .A(B[4]), .Y(n998) );
  INVX2 U1383 ( .A(n1000), .Y(n1001) );
  INVX2 U1384 ( .A(B[5]), .Y(n1000) );
  INVX1 U1385 ( .A(n984), .Y(n1044) );
  INVX1 U1386 ( .A(n985), .Y(n1043) );
  INVX4 U1387 ( .A(B[2]), .Y(n994) );
  INVX8 U1388 ( .A(n990), .Y(n991) );
  INVX8 U1389 ( .A(n994), .Y(n995) );
  INVX8 U1390 ( .A(n1008), .Y(n1009) );
  INVX8 U1391 ( .A(n1012), .Y(n1013) );
  INVX8 U1392 ( .A(n1014), .Y(n1015) );
  INVX8 U1393 ( .A(n1016), .Y(n1017) );
  INVX8 U1394 ( .A(n1018), .Y(n1019) );
  INVX8 U1395 ( .A(n1024), .Y(n1025) );
  INVX8 U1396 ( .A(n1026), .Y(n1027) );
  INVX8 U1397 ( .A(n1028), .Y(n1029) );
  INVX8 U1398 ( .A(n1030), .Y(n1031) );
  INVX8 U1399 ( .A(n1032), .Y(n1033) );
  INVX8 U1400 ( .A(n1034), .Y(n1035) );
  INVX8 U1401 ( .A(n1036), .Y(n1037) );
  AND2X2 U1402 ( .A(n846), .B(n1019), .Y(\ab[1][14] ) );
  AND2X2 U1403 ( .A(n1019), .B(n987), .Y(\ab[0][14] ) );
  AND2X2 U1404 ( .A(n322), .B(n1017), .Y(\ab[1][13] ) );
  AND2X2 U1405 ( .A(n1017), .B(n266), .Y(\ab[0][13] ) );
  AND2X2 U1406 ( .A(n511), .B(n1015), .Y(\ab[1][12] ) );
  AND2X2 U1407 ( .A(n322), .B(n1013), .Y(\ab[1][11] ) );
  AND2X2 U1408 ( .A(n1013), .B(n987), .Y(\ab[0][11] ) );
  AND2X2 U1409 ( .A(n511), .B(B[10]), .Y(\ab[1][10] ) );
  AND2X2 U1410 ( .A(n266), .B(B[10]), .Y(\ab[0][10] ) );
  AND2X2 U1411 ( .A(n266), .B(B[9]), .Y(\ab[0][9] ) );
  AND2X2 U1412 ( .A(n1007), .B(n514), .Y(\ab[1][8] ) );
  AND2X2 U1413 ( .A(n266), .B(n239), .Y(\ab[0][8] ) );
  AND2X2 U1414 ( .A(B[7]), .B(n987), .Y(\ab[0][7] ) );
  AND2X2 U1415 ( .A(B[6]), .B(n514), .Y(\ab[1][6] ) );
  AND2X2 U1416 ( .A(n1001), .B(n514), .Y(\ab[1][5] ) );
  AND2X2 U1417 ( .A(n1001), .B(n266), .Y(\ab[0][5] ) );
  AND2X2 U1418 ( .A(n999), .B(n987), .Y(\ab[0][4] ) );
  AND2X2 U1419 ( .A(n997), .B(n514), .Y(\ab[1][3] ) );
  AND2X2 U1420 ( .A(n997), .B(n987), .Y(\ab[0][3] ) );
  AND2X2 U1421 ( .A(n995), .B(n987), .Y(\ab[0][2] ) );
  AND2X2 U1422 ( .A(n993), .B(n987), .Y(\ab[0][1] ) );
  AND2X2 U1423 ( .A(n991), .B(n846), .Y(\ab[1][0] ) );
  AND2X2 U1424 ( .A(n235), .B(n1019), .Y(\ab[2][14] ) );
  NOR2X1 U1425 ( .A(n846), .B(n1049), .Y(\ab[1][15] ) );
  AND2X2 U1426 ( .A(n236), .B(n1017), .Y(\ab[2][13] ) );
  AND2X2 U1427 ( .A(n235), .B(n1015), .Y(\ab[2][12] ) );
  AND2X2 U1428 ( .A(n236), .B(n1013), .Y(\ab[2][11] ) );
  AND2X2 U1429 ( .A(n235), .B(n51), .Y(\ab[2][10] ) );
  AND2X2 U1430 ( .A(n206), .B(B[9]), .Y(\ab[2][9] ) );
  AND2X2 U1431 ( .A(n1023), .B(B[6]), .Y(\ab[2][6] ) );
  AND2X2 U1432 ( .A(n236), .B(n983), .Y(\ab[2][3] ) );
  AND2X2 U1433 ( .A(n1023), .B(n995), .Y(\ab[2][2] ) );
  AND2X2 U1434 ( .A(n235), .B(n991), .Y(\ab[2][0] ) );
  AND2X2 U1435 ( .A(n1025), .B(n1019), .Y(\ab[3][14] ) );
  NOR2X1 U1436 ( .A(n235), .B(n1049), .Y(\ab[2][15] ) );
  AND2X2 U1437 ( .A(n1025), .B(n1017), .Y(\ab[3][13] ) );
  AND2X2 U1438 ( .A(n1025), .B(n1015), .Y(\ab[3][12] ) );
  AND2X2 U1439 ( .A(n1025), .B(n1013), .Y(\ab[3][11] ) );
  AND2X2 U1440 ( .A(n1025), .B(n51), .Y(\ab[3][10] ) );
  AND2X2 U1441 ( .A(n1025), .B(B[7]), .Y(\ab[3][7] ) );
  AND2X2 U1442 ( .A(n1025), .B(n1003), .Y(\ab[3][6] ) );
  AND2X2 U1443 ( .A(n1025), .B(n985), .Y(\ab[3][5] ) );
  AND2X2 U1444 ( .A(n1025), .B(n984), .Y(\ab[3][4] ) );
  AND2X2 U1445 ( .A(n1025), .B(n983), .Y(\ab[3][3] ) );
  AND2X2 U1446 ( .A(n1025), .B(n995), .Y(\ab[3][2] ) );
  AND2X2 U1447 ( .A(n1025), .B(n993), .Y(\ab[3][1] ) );
  AND2X2 U1448 ( .A(n396), .B(n991), .Y(\ab[3][0] ) );
  AND2X2 U1449 ( .A(n1027), .B(n1019), .Y(\ab[4][14] ) );
  NOR2X1 U1450 ( .A(n396), .B(n1049), .Y(\ab[3][15] ) );
  AND2X2 U1451 ( .A(n1027), .B(n1017), .Y(\ab[4][13] ) );
  AND2X2 U1452 ( .A(n1027), .B(n1015), .Y(\ab[4][12] ) );
  AND2X2 U1453 ( .A(n1027), .B(n1013), .Y(\ab[4][11] ) );
  AND2X2 U1454 ( .A(n1027), .B(n1011), .Y(\ab[4][10] ) );
  AND2X2 U1455 ( .A(n1027), .B(n1009), .Y(\ab[4][9] ) );
  AND2X2 U1456 ( .A(n1027), .B(n1007), .Y(\ab[4][8] ) );
  AND2X2 U1457 ( .A(n1027), .B(n1005), .Y(\ab[4][7] ) );
  AND2X2 U1458 ( .A(n1027), .B(n1003), .Y(\ab[4][6] ) );
  AND2X2 U1459 ( .A(n1027), .B(n985), .Y(\ab[4][5] ) );
  AND2X2 U1460 ( .A(n1027), .B(n984), .Y(\ab[4][4] ) );
  AND2X2 U1461 ( .A(n1027), .B(n983), .Y(\ab[4][3] ) );
  AND2X2 U1462 ( .A(n1027), .B(n995), .Y(\ab[4][2] ) );
  AND2X2 U1463 ( .A(n1027), .B(n993), .Y(\ab[4][1] ) );
  AND2X2 U1464 ( .A(n1027), .B(n991), .Y(\ab[4][0] ) );
  AND2X2 U1465 ( .A(n1029), .B(n1019), .Y(\ab[5][14] ) );
  NOR2X1 U1466 ( .A(n1027), .B(n1049), .Y(\ab[4][15] ) );
  AND2X2 U1467 ( .A(n1029), .B(n1017), .Y(\ab[5][13] ) );
  AND2X2 U1468 ( .A(n1029), .B(n1015), .Y(\ab[5][12] ) );
  AND2X2 U1469 ( .A(n1029), .B(n1013), .Y(\ab[5][11] ) );
  AND2X2 U1470 ( .A(n1029), .B(n1011), .Y(\ab[5][10] ) );
  AND2X2 U1471 ( .A(n1029), .B(n1009), .Y(\ab[5][9] ) );
  AND2X2 U1472 ( .A(n1029), .B(n1007), .Y(\ab[5][8] ) );
  AND2X2 U1473 ( .A(n1029), .B(n1005), .Y(\ab[5][7] ) );
  AND2X2 U1474 ( .A(n1029), .B(n1003), .Y(\ab[5][6] ) );
  AND2X2 U1475 ( .A(n1029), .B(n985), .Y(\ab[5][5] ) );
  AND2X2 U1476 ( .A(n1029), .B(n984), .Y(\ab[5][4] ) );
  AND2X2 U1477 ( .A(n1029), .B(n983), .Y(\ab[5][3] ) );
  AND2X2 U1478 ( .A(n1029), .B(n995), .Y(\ab[5][2] ) );
  AND2X2 U1479 ( .A(n1029), .B(n993), .Y(\ab[5][1] ) );
  AND2X2 U1480 ( .A(n1029), .B(n991), .Y(\ab[5][0] ) );
  AND2X2 U1481 ( .A(n1031), .B(n1019), .Y(\ab[6][14] ) );
  NOR2X1 U1482 ( .A(n1029), .B(n1049), .Y(\ab[5][15] ) );
  AND2X2 U1483 ( .A(n1031), .B(n1017), .Y(\ab[6][13] ) );
  AND2X2 U1484 ( .A(n1031), .B(n1015), .Y(\ab[6][12] ) );
  AND2X2 U1485 ( .A(n1031), .B(n1013), .Y(\ab[6][11] ) );
  AND2X2 U1486 ( .A(n1031), .B(n1011), .Y(\ab[6][10] ) );
  AND2X2 U1487 ( .A(n1031), .B(n1009), .Y(\ab[6][9] ) );
  AND2X2 U1488 ( .A(n1031), .B(n1007), .Y(\ab[6][8] ) );
  AND2X2 U1489 ( .A(n1031), .B(n1005), .Y(\ab[6][7] ) );
  AND2X2 U1490 ( .A(n1031), .B(n1003), .Y(\ab[6][6] ) );
  AND2X2 U1491 ( .A(n1031), .B(n985), .Y(\ab[6][5] ) );
  AND2X2 U1492 ( .A(n1031), .B(n984), .Y(\ab[6][4] ) );
  AND2X2 U1493 ( .A(n1031), .B(n983), .Y(\ab[6][3] ) );
  AND2X2 U1494 ( .A(n1031), .B(n995), .Y(\ab[6][2] ) );
  AND2X2 U1495 ( .A(n1031), .B(n993), .Y(\ab[6][1] ) );
  AND2X2 U1496 ( .A(n1031), .B(n991), .Y(\ab[6][0] ) );
  AND2X2 U1497 ( .A(n1033), .B(n1019), .Y(\ab[7][14] ) );
  NOR2X1 U1498 ( .A(n1031), .B(n1049), .Y(\ab[6][15] ) );
  AND2X2 U1499 ( .A(n1033), .B(n1017), .Y(\ab[7][13] ) );
  AND2X2 U1500 ( .A(n1033), .B(n1015), .Y(\ab[7][12] ) );
  AND2X2 U1501 ( .A(n1033), .B(n1013), .Y(\ab[7][11] ) );
  AND2X2 U1502 ( .A(n1033), .B(n1011), .Y(\ab[7][10] ) );
  AND2X2 U1503 ( .A(n1033), .B(n1009), .Y(\ab[7][9] ) );
  AND2X2 U1504 ( .A(n1033), .B(n132), .Y(\ab[7][8] ) );
  AND2X2 U1505 ( .A(n1033), .B(n1005), .Y(\ab[7][7] ) );
  AND2X2 U1506 ( .A(n1033), .B(n1003), .Y(\ab[7][6] ) );
  AND2X2 U1507 ( .A(n1033), .B(n985), .Y(\ab[7][5] ) );
  AND2X2 U1508 ( .A(n1033), .B(n984), .Y(\ab[7][4] ) );
  AND2X2 U1509 ( .A(n1033), .B(n983), .Y(\ab[7][3] ) );
  AND2X2 U1510 ( .A(n1033), .B(n995), .Y(\ab[7][2] ) );
  AND2X2 U1511 ( .A(n1033), .B(n993), .Y(\ab[7][1] ) );
  AND2X2 U1512 ( .A(n1033), .B(n991), .Y(\ab[7][0] ) );
  AND2X2 U1513 ( .A(n1035), .B(n1019), .Y(\ab[8][14] ) );
  NOR2X1 U1514 ( .A(n1033), .B(n1049), .Y(\ab[7][15] ) );
  AND2X2 U1515 ( .A(n1035), .B(n1017), .Y(\ab[8][13] ) );
  AND2X2 U1516 ( .A(n1035), .B(n1015), .Y(\ab[8][12] ) );
  AND2X2 U1517 ( .A(n1035), .B(n1013), .Y(\ab[8][11] ) );
  AND2X2 U1518 ( .A(n1035), .B(n1011), .Y(\ab[8][10] ) );
  AND2X2 U1519 ( .A(n1035), .B(n1009), .Y(\ab[8][9] ) );
  AND2X2 U1520 ( .A(n1035), .B(n132), .Y(\ab[8][8] ) );
  AND2X2 U1521 ( .A(n1035), .B(n1005), .Y(\ab[8][7] ) );
  AND2X2 U1522 ( .A(n1035), .B(n1003), .Y(\ab[8][6] ) );
  AND2X2 U1523 ( .A(n1035), .B(n985), .Y(\ab[8][5] ) );
  AND2X2 U1524 ( .A(n1035), .B(n984), .Y(\ab[8][4] ) );
  AND2X2 U1525 ( .A(n1035), .B(n983), .Y(\ab[8][3] ) );
  AND2X2 U1526 ( .A(n1035), .B(n995), .Y(\ab[8][2] ) );
  AND2X2 U1527 ( .A(n1035), .B(n993), .Y(\ab[8][1] ) );
  AND2X2 U1528 ( .A(n1035), .B(n991), .Y(\ab[8][0] ) );
  AND2X2 U1529 ( .A(n1037), .B(n1019), .Y(\ab[9][14] ) );
  NOR2X1 U1530 ( .A(n1035), .B(n1049), .Y(\ab[8][15] ) );
  AND2X2 U1531 ( .A(n1037), .B(n1017), .Y(\ab[9][13] ) );
  AND2X2 U1532 ( .A(n1037), .B(n1015), .Y(\ab[9][12] ) );
  AND2X2 U1533 ( .A(n1037), .B(n1013), .Y(\ab[9][11] ) );
  AND2X2 U1534 ( .A(n1037), .B(n1011), .Y(\ab[9][10] ) );
  AND2X2 U1535 ( .A(n1037), .B(n1009), .Y(\ab[9][9] ) );
  AND2X2 U1536 ( .A(n1037), .B(n132), .Y(\ab[9][8] ) );
  AND2X2 U1537 ( .A(n1037), .B(n1005), .Y(\ab[9][7] ) );
  AND2X2 U1538 ( .A(n1037), .B(n1003), .Y(\ab[9][6] ) );
  AND2X2 U1539 ( .A(n1037), .B(n985), .Y(\ab[9][5] ) );
  AND2X2 U1540 ( .A(n1037), .B(n984), .Y(\ab[9][4] ) );
  AND2X2 U1541 ( .A(n1037), .B(n983), .Y(\ab[9][3] ) );
  AND2X2 U1542 ( .A(n1037), .B(n995), .Y(\ab[9][2] ) );
  AND2X2 U1543 ( .A(n1037), .B(n993), .Y(\ab[9][1] ) );
  AND2X2 U1544 ( .A(n1037), .B(n991), .Y(\ab[9][0] ) );
  AND2X2 U1545 ( .A(A[10]), .B(n1019), .Y(\ab[10][14] ) );
  NOR2X1 U1546 ( .A(n1037), .B(n1049), .Y(\ab[9][15] ) );
  AND2X2 U1547 ( .A(A[10]), .B(n1017), .Y(\ab[10][13] ) );
  AND2X2 U1548 ( .A(A[10]), .B(n1015), .Y(\ab[10][12] ) );
  AND2X2 U1549 ( .A(A[10]), .B(n1013), .Y(\ab[10][11] ) );
  AND2X2 U1550 ( .A(A[10]), .B(n1011), .Y(\ab[10][10] ) );
  AND2X2 U1551 ( .A(A[10]), .B(n1009), .Y(\ab[10][9] ) );
  AND2X2 U1552 ( .A(A[10]), .B(n132), .Y(\ab[10][8] ) );
  AND2X2 U1553 ( .A(A[10]), .B(n1005), .Y(\ab[10][7] ) );
  AND2X2 U1554 ( .A(A[10]), .B(n1003), .Y(\ab[10][6] ) );
  AND2X2 U1555 ( .A(A[10]), .B(n985), .Y(\ab[10][5] ) );
  AND2X2 U1556 ( .A(A[10]), .B(n984), .Y(\ab[10][4] ) );
  AND2X2 U1557 ( .A(A[10]), .B(n983), .Y(\ab[10][3] ) );
  AND2X2 U1558 ( .A(A[10]), .B(n995), .Y(\ab[10][2] ) );
  AND2X2 U1559 ( .A(A[10]), .B(n993), .Y(\ab[10][1] ) );
  AND2X2 U1560 ( .A(A[10]), .B(n991), .Y(\ab[10][0] ) );
  AND2X2 U1561 ( .A(A[11]), .B(n1019), .Y(\ab[11][14] ) );
  NOR2X1 U1562 ( .A(A[10]), .B(n1049), .Y(\ab[10][15] ) );
  AND2X2 U1563 ( .A(A[11]), .B(n1017), .Y(\ab[11][13] ) );
  AND2X2 U1564 ( .A(A[11]), .B(n1015), .Y(\ab[11][12] ) );
  AND2X2 U1565 ( .A(A[11]), .B(n1013), .Y(\ab[11][11] ) );
  AND2X2 U1566 ( .A(A[11]), .B(n1011), .Y(\ab[11][10] ) );
  AND2X2 U1567 ( .A(A[11]), .B(n1009), .Y(\ab[11][9] ) );
  AND2X2 U1568 ( .A(A[11]), .B(n132), .Y(\ab[11][8] ) );
  AND2X2 U1569 ( .A(A[11]), .B(n1005), .Y(\ab[11][7] ) );
  AND2X2 U1570 ( .A(A[11]), .B(n1003), .Y(\ab[11][6] ) );
  AND2X2 U1571 ( .A(A[11]), .B(n985), .Y(\ab[11][5] ) );
  AND2X2 U1572 ( .A(A[11]), .B(n984), .Y(\ab[11][4] ) );
  AND2X2 U1573 ( .A(A[11]), .B(n983), .Y(\ab[11][3] ) );
  AND2X2 U1574 ( .A(A[11]), .B(n995), .Y(\ab[11][2] ) );
  AND2X2 U1575 ( .A(A[11]), .B(n993), .Y(\ab[11][1] ) );
  AND2X2 U1576 ( .A(A[11]), .B(n991), .Y(\ab[11][0] ) );
  AND2X2 U1577 ( .A(A[12]), .B(n1019), .Y(\ab[12][14] ) );
  NOR2X1 U1578 ( .A(A[11]), .B(n1049), .Y(\ab[11][15] ) );
  AND2X2 U1579 ( .A(A[12]), .B(n1017), .Y(\ab[12][13] ) );
  AND2X2 U1580 ( .A(A[12]), .B(n1015), .Y(\ab[12][12] ) );
  AND2X2 U1581 ( .A(A[12]), .B(n1013), .Y(\ab[12][11] ) );
  AND2X2 U1582 ( .A(A[12]), .B(n1011), .Y(\ab[12][10] ) );
  AND2X2 U1583 ( .A(A[12]), .B(n1009), .Y(\ab[12][9] ) );
  AND2X2 U1584 ( .A(A[12]), .B(n132), .Y(\ab[12][8] ) );
  AND2X2 U1585 ( .A(A[12]), .B(n1005), .Y(\ab[12][7] ) );
  AND2X2 U1586 ( .A(A[12]), .B(n1003), .Y(\ab[12][6] ) );
  AND2X2 U1587 ( .A(A[12]), .B(n985), .Y(\ab[12][5] ) );
  AND2X2 U1588 ( .A(A[12]), .B(n984), .Y(\ab[12][4] ) );
  AND2X2 U1589 ( .A(A[12]), .B(n983), .Y(\ab[12][3] ) );
  AND2X2 U1590 ( .A(A[12]), .B(n995), .Y(\ab[12][2] ) );
  AND2X2 U1591 ( .A(A[12]), .B(n993), .Y(\ab[12][1] ) );
  AND2X2 U1592 ( .A(A[12]), .B(n991), .Y(\ab[12][0] ) );
  NOR2X1 U1593 ( .A(n1052), .B(n1018), .Y(\ab[13][14] ) );
  NOR2X1 U1594 ( .A(A[12]), .B(n1049), .Y(\ab[12][15] ) );
  NOR2X1 U1595 ( .A(n1052), .B(n1038), .Y(\ab[13][13] ) );
  NOR2X1 U1596 ( .A(n1052), .B(n1039), .Y(\ab[13][12] ) );
  NOR2X1 U1597 ( .A(n1052), .B(n1040), .Y(\ab[13][11] ) );
  NOR2X1 U1598 ( .A(n1052), .B(n1010), .Y(\ab[13][10] ) );
  NOR2X1 U1599 ( .A(n1052), .B(n1041), .Y(\ab[13][9] ) );
  NOR2X1 U1600 ( .A(n1052), .B(n1042), .Y(\ab[13][8] ) );
  NOR2X1 U1601 ( .A(n1052), .B(n1004), .Y(\ab[13][7] ) );
  NOR2X1 U1602 ( .A(n1052), .B(n1002), .Y(\ab[13][6] ) );
  NOR2X1 U1603 ( .A(n1052), .B(n1043), .Y(\ab[13][5] ) );
  NOR2X1 U1604 ( .A(n1052), .B(n1044), .Y(\ab[13][4] ) );
  NOR2X1 U1605 ( .A(n1052), .B(n996), .Y(\ab[13][3] ) );
  INVX2 U1606 ( .A(n995), .Y(n1045) );
  NOR2X1 U1607 ( .A(n1052), .B(n1045), .Y(\ab[13][2] ) );
  INVX2 U1608 ( .A(n993), .Y(n1046) );
  NOR2X1 U1609 ( .A(n1052), .B(n1046), .Y(\ab[13][1] ) );
  INVX2 U1610 ( .A(n991), .Y(n1047) );
  NOR2X1 U1611 ( .A(n1052), .B(n1047), .Y(\ab[13][0] ) );
  NOR2X1 U1612 ( .A(n1051), .B(n1018), .Y(\ab[14][14] ) );
  NOR2X1 U1613 ( .A(A[13]), .B(n1049), .Y(\ab[13][15] ) );
  NOR2X1 U1614 ( .A(n1051), .B(n1038), .Y(\ab[14][13] ) );
  NOR2X1 U1615 ( .A(n1051), .B(n1039), .Y(\ab[14][12] ) );
  NOR2X1 U1616 ( .A(n1051), .B(n1040), .Y(\ab[14][11] ) );
  NOR2X1 U1617 ( .A(n1051), .B(n1010), .Y(\ab[14][10] ) );
  NOR2X1 U1618 ( .A(n1051), .B(n1041), .Y(\ab[14][9] ) );
  NOR2X1 U1619 ( .A(n1051), .B(n1042), .Y(\ab[14][8] ) );
  NOR2X1 U1620 ( .A(n1051), .B(n1004), .Y(\ab[14][7] ) );
  NOR2X1 U1621 ( .A(n1051), .B(n1002), .Y(\ab[14][6] ) );
  NOR2X1 U1622 ( .A(n1051), .B(n1043), .Y(\ab[14][5] ) );
  NOR2X1 U1623 ( .A(n1051), .B(n1044), .Y(\ab[14][4] ) );
  NOR2X1 U1624 ( .A(n1051), .B(n996), .Y(\ab[14][3] ) );
  NOR2X1 U1625 ( .A(n1051), .B(n1045), .Y(\ab[14][2] ) );
  NOR2X1 U1626 ( .A(n1051), .B(n1046), .Y(\ab[14][1] ) );
  NOR2X1 U1627 ( .A(n1051), .B(n1047), .Y(\ab[14][0] ) );
  NOR2X1 U1628 ( .A(n1050), .B(n1049), .Y(\ab[15][15] ) );
  NOR2X1 U1629 ( .A(A[14]), .B(n1049), .Y(\ab[14][15] ) );
  AND2X2 U1630 ( .A(n991), .B(n987), .Y(PRODUCT[0]) );
  INVX2 U1631 ( .A(\CARRYB[15][15] ), .Y(n1048) );
  NOR2X1 U1632 ( .A(n1009), .B(n1050), .Y(\ab[15][9] ) );
  NOR2X1 U1633 ( .A(n132), .B(n1050), .Y(\ab[15][8] ) );
  NOR2X1 U1634 ( .A(n1005), .B(n1050), .Y(\ab[15][7] ) );
  NOR2X1 U1635 ( .A(n1003), .B(n1050), .Y(\ab[15][6] ) );
  NOR2X1 U1636 ( .A(n985), .B(n1050), .Y(\ab[15][5] ) );
  NOR2X1 U1637 ( .A(n984), .B(n1050), .Y(\ab[15][4] ) );
  NOR2X1 U1638 ( .A(n983), .B(n1050), .Y(\ab[15][3] ) );
  NOR2X1 U1639 ( .A(n995), .B(n1050), .Y(\ab[15][2] ) );
  NOR2X1 U1640 ( .A(n993), .B(n1050), .Y(\ab[15][1] ) );
  NOR2X1 U1641 ( .A(n1019), .B(n1050), .Y(\ab[15][14] ) );
  NOR2X1 U1642 ( .A(n1017), .B(n1050), .Y(\ab[15][13] ) );
  NOR2X1 U1643 ( .A(n1015), .B(n1050), .Y(\ab[15][12] ) );
  NOR2X1 U1644 ( .A(n1013), .B(n1050), .Y(\ab[15][11] ) );
  NOR2X1 U1645 ( .A(n1011), .B(n1050), .Y(\ab[15][10] ) );
  NOR2X1 U1646 ( .A(n991), .B(n1050), .Y(\ab[15][0] ) );
endmodule


module matrix_math_DW01_add_13 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160;

  NAND3X1 U2 ( .A(n74), .B(n73), .C(n72), .Y(n1) );
  OR2X1 U3 ( .A(A[22]), .B(B[22]), .Y(n66) );
  AND2X2 U4 ( .A(A[22]), .B(B[22]), .Y(n6) );
  XNOR2X1 U5 ( .A(n13), .B(n2), .Y(SUM[21]) );
  NAND2X1 U6 ( .A(n79), .B(n72), .Y(n2) );
  NAND2X1 U7 ( .A(n3), .B(n4), .Y(n5) );
  NAND2X1 U8 ( .A(n5), .B(n101), .Y(n100) );
  INVX1 U9 ( .A(n19), .Y(n3) );
  INVX2 U10 ( .A(n98), .Y(n4) );
  AND2X2 U11 ( .A(n87), .B(n86), .Y(SUM[0]) );
  XNOR2X1 U12 ( .A(A[22]), .B(B[22]), .Y(n67) );
  AND2X1 U13 ( .A(n103), .B(n10), .Y(n101) );
  NOR2X1 U14 ( .A(B[17]), .B(A[17]), .Y(n8) );
  INVX2 U15 ( .A(n26), .Y(n27) );
  OAI21X1 U16 ( .A(n69), .B(n70), .C(n71), .Y(n9) );
  OR2X2 U17 ( .A(B[17]), .B(A[17]), .Y(n10) );
  BUFX2 U18 ( .A(A[18]), .Y(n11) );
  XOR2X1 U19 ( .A(n64), .B(n12), .Y(SUM[23]) );
  XNOR2X1 U20 ( .A(B[23]), .B(A[23]), .Y(n12) );
  NAND2X1 U21 ( .A(n71), .B(n74), .Y(n13) );
  XOR2X1 U22 ( .A(n99), .B(n14), .Y(SUM[18]) );
  AND2X2 U23 ( .A(n94), .B(n93), .Y(n14) );
  XOR2X1 U24 ( .A(n67), .B(n9), .Y(SUM[22]) );
  NOR2X1 U25 ( .A(n15), .B(n8), .Y(n90) );
  INVX1 U26 ( .A(n15), .Y(n94) );
  NOR2X1 U27 ( .A(A[18]), .B(B[18]), .Y(n15) );
  AND2X2 U28 ( .A(B[16]), .B(A[16]), .Y(n19) );
  INVX1 U29 ( .A(n137), .Y(n147) );
  INVX1 U30 ( .A(n42), .Y(n41) );
  XOR2X1 U31 ( .A(n83), .B(n84), .Y(SUM[20]) );
  XOR2X1 U32 ( .A(n27), .B(n88), .Y(SUM[19]) );
  XOR2X1 U33 ( .A(n102), .B(n17), .Y(SUM[17]) );
  NAND2X1 U34 ( .A(n10), .B(n92), .Y(n17) );
  XNOR2X1 U35 ( .A(n124), .B(n125), .Y(SUM[15]) );
  XNOR2X1 U36 ( .A(n127), .B(n18), .Y(SUM[14]) );
  NAND2X1 U37 ( .A(n107), .B(n112), .Y(n18) );
  XOR2X1 U38 ( .A(n104), .B(n98), .Y(SUM[16]) );
  XOR2X1 U39 ( .A(n133), .B(n20), .Y(SUM[12]) );
  NAND2X1 U40 ( .A(n122), .B(n117), .Y(n20) );
  XOR2X1 U41 ( .A(n144), .B(n145), .Y(SUM[11]) );
  NOR2X1 U42 ( .A(n142), .B(n143), .Y(n21) );
  XNOR2X1 U43 ( .A(n146), .B(n22), .Y(SUM[10]) );
  NAND2X1 U44 ( .A(n141), .B(n137), .Y(n22) );
  XOR2X1 U45 ( .A(n28), .B(n23), .Y(SUM[9]) );
  NAND2X1 U46 ( .A(n29), .B(n30), .Y(n23) );
  XNOR2X1 U47 ( .A(n39), .B(n24), .Y(SUM[6]) );
  NAND2X1 U48 ( .A(n40), .B(n42), .Y(n24) );
  XNOR2X1 U49 ( .A(n31), .B(n32), .Y(SUM[8]) );
  XOR2X1 U50 ( .A(n35), .B(n36), .Y(SUM[7]) );
  XNOR2X1 U51 ( .A(n45), .B(n25), .Y(SUM[5]) );
  NAND2X1 U52 ( .A(n46), .B(n44), .Y(n25) );
  INVX2 U53 ( .A(n86), .Y(n62) );
  NAND2X1 U54 ( .A(n115), .B(n116), .Y(n114) );
  INVX2 U55 ( .A(n81), .Y(n26) );
  NAND2X1 U56 ( .A(n33), .B(n34), .Y(n32) );
  NAND2X1 U57 ( .A(n37), .B(n38), .Y(n36) );
  AOI21X1 U58 ( .A(n39), .B(n40), .C(n41), .Y(n35) );
  NAND2X1 U59 ( .A(n43), .B(n44), .Y(n39) );
  NAND2X1 U60 ( .A(n45), .B(n46), .Y(n43) );
  OAI21X1 U61 ( .A(n119), .B(n47), .C(n48), .Y(n45) );
  INVX2 U62 ( .A(n49), .Y(n47) );
  XNOR2X1 U63 ( .A(n50), .B(n155), .Y(SUM[4]) );
  NAND2X1 U64 ( .A(n48), .B(n49), .Y(n50) );
  XNOR2X1 U65 ( .A(n51), .B(n52), .Y(SUM[3]) );
  AND2X2 U66 ( .A(n53), .B(n54), .Y(n52) );
  AOI21X1 U67 ( .A(n55), .B(n56), .C(n57), .Y(n51) );
  INVX2 U68 ( .A(n58), .Y(n57) );
  XNOR2X1 U69 ( .A(n59), .B(n60), .Y(SUM[2]) );
  AND2X2 U70 ( .A(n56), .B(n58), .Y(n60) );
  INVX2 U71 ( .A(n55), .Y(n59) );
  OAI21X1 U72 ( .A(n160), .B(n86), .C(n61), .Y(n55) );
  AOI21X1 U73 ( .A(n66), .B(n65), .C(n6), .Y(n64) );
  INVX2 U74 ( .A(n68), .Y(n65) );
  OAI21X1 U75 ( .A(n69), .B(n1), .C(n71), .Y(n68) );
  NAND3X1 U76 ( .A(n74), .B(n73), .C(n72), .Y(n70) );
  NAND2X1 U77 ( .A(n76), .B(n75), .Y(n73) );
  INVX2 U78 ( .A(n77), .Y(n69) );
  NAND3X1 U79 ( .A(n78), .B(n76), .C(n26), .Y(n77) );
  NAND2X1 U80 ( .A(B[21]), .B(A[21]), .Y(n74) );
  OR2X2 U81 ( .A(A[21]), .B(B[21]), .Y(n71) );
  NAND3X1 U82 ( .A(n78), .B(n76), .C(n80), .Y(n79) );
  NAND2X1 U83 ( .A(n82), .B(n81), .Y(n80) );
  NAND2X1 U84 ( .A(n72), .B(n76), .Y(n84) );
  OR2X2 U85 ( .A(A[20]), .B(B[20]), .Y(n76) );
  NAND2X1 U86 ( .A(B[20]), .B(A[20]), .Y(n72) );
  AOI21X1 U87 ( .A(n26), .B(n78), .C(n75), .Y(n83) );
  INVX2 U88 ( .A(n82), .Y(n75) );
  XNOR2X1 U89 ( .A(n85), .B(n62), .Y(SUM[1]) );
  NAND2X1 U90 ( .A(n63), .B(n61), .Y(n85) );
  AOI21X1 U91 ( .A(n89), .B(n90), .C(n91), .Y(n81) );
  OAI21X1 U92 ( .A(n15), .B(n92), .C(n93), .Y(n91) );
  AOI21X1 U93 ( .A(n95), .B(n96), .C(n97), .Y(n89) );
  NOR2X1 U94 ( .A(B[16]), .B(A[16]), .Y(n97) );
  INVX2 U95 ( .A(n98), .Y(n96) );
  NAND2X1 U96 ( .A(B[16]), .B(A[16]), .Y(n95) );
  NAND2X1 U97 ( .A(n82), .B(n78), .Y(n88) );
  OR2X2 U98 ( .A(B[19]), .B(A[19]), .Y(n78) );
  NAND2X1 U99 ( .A(B[19]), .B(A[19]), .Y(n82) );
  NAND2X1 U100 ( .A(n11), .B(B[18]), .Y(n93) );
  NAND2X1 U101 ( .A(n92), .B(n100), .Y(n99) );
  NAND2X1 U102 ( .A(B[17]), .B(A[17]), .Y(n92) );
  AOI21X1 U103 ( .A(n98), .B(n103), .C(n19), .Y(n102) );
  OR2X2 U104 ( .A(A[16]), .B(B[16]), .Y(n103) );
  NAND2X1 U105 ( .A(n105), .B(n106), .Y(n98) );
  NAND3X1 U106 ( .A(n107), .B(n108), .C(n109), .Y(n106) );
  NAND3X1 U107 ( .A(n110), .B(n111), .C(n112), .Y(n108) );
  NAND2X1 U108 ( .A(n113), .B(n114), .Y(n111) );
  AND2X2 U109 ( .A(n117), .B(n118), .Y(n116) );
  NAND2X1 U110 ( .A(n21), .B(n31), .Y(n115) );
  AND2X2 U111 ( .A(n122), .B(n123), .Y(n113) );
  XOR2X1 U112 ( .A(B[16]), .B(A[16]), .Y(n104) );
  NAND2X1 U113 ( .A(n105), .B(n109), .Y(n125) );
  OR2X2 U114 ( .A(A[15]), .B(B[15]), .Y(n109) );
  NAND2X1 U115 ( .A(B[15]), .B(A[15]), .Y(n105) );
  NAND2X1 U116 ( .A(n112), .B(n126), .Y(n124) );
  NAND2X1 U117 ( .A(n127), .B(n107), .Y(n126) );
  NAND2X1 U118 ( .A(B[14]), .B(A[14]), .Y(n112) );
  OR2X2 U119 ( .A(A[14]), .B(B[14]), .Y(n107) );
  OAI21X1 U120 ( .A(n128), .B(n129), .C(n110), .Y(n127) );
  INVX2 U121 ( .A(n130), .Y(n129) );
  INVX2 U122 ( .A(n123), .Y(n128) );
  XNOR2X1 U123 ( .A(n131), .B(n130), .Y(SUM[13]) );
  OAI21X1 U124 ( .A(n132), .B(n133), .C(n117), .Y(n130) );
  INVX2 U125 ( .A(n122), .Y(n132) );
  NAND2X1 U126 ( .A(n123), .B(n110), .Y(n131) );
  NAND2X1 U127 ( .A(B[13]), .B(A[13]), .Y(n110) );
  OR2X2 U128 ( .A(A[13]), .B(B[13]), .Y(n123) );
  NAND2X1 U129 ( .A(B[12]), .B(A[12]), .Y(n117) );
  OR2X2 U130 ( .A(A[12]), .B(B[12]), .Y(n122) );
  AND2X2 U131 ( .A(n134), .B(n118), .Y(n133) );
  NAND2X1 U132 ( .A(n135), .B(n136), .Y(n118) );
  NAND3X1 U133 ( .A(n137), .B(n138), .C(n139), .Y(n136) );
  NAND3X1 U134 ( .A(n29), .B(n140), .C(n141), .Y(n138) );
  NAND2X1 U135 ( .A(n30), .B(n33), .Y(n140) );
  NAND2X1 U136 ( .A(n21), .B(n31), .Y(n134) );
  NAND3X1 U137 ( .A(n29), .B(n34), .C(n141), .Y(n143) );
  INVX2 U138 ( .A(n135), .Y(n142) );
  NAND2X1 U139 ( .A(n139), .B(n135), .Y(n145) );
  OR2X2 U140 ( .A(A[11]), .B(B[11]), .Y(n135) );
  NAND2X1 U141 ( .A(B[11]), .B(A[11]), .Y(n139) );
  AOI21X1 U142 ( .A(n146), .B(n141), .C(n147), .Y(n144) );
  NAND2X1 U143 ( .A(B[10]), .B(A[10]), .Y(n137) );
  OR2X2 U144 ( .A(A[10]), .B(B[10]), .Y(n141) );
  OAI21X1 U145 ( .A(n28), .B(n148), .C(n30), .Y(n146) );
  NAND2X1 U146 ( .A(B[9]), .B(A[9]), .Y(n30) );
  INVX2 U147 ( .A(n29), .Y(n148) );
  OR2X2 U148 ( .A(A[9]), .B(B[9]), .Y(n29) );
  AND2X2 U149 ( .A(n149), .B(n33), .Y(n28) );
  NAND2X1 U150 ( .A(B[8]), .B(A[8]), .Y(n33) );
  NAND2X1 U151 ( .A(n34), .B(n31), .Y(n149) );
  OAI21X1 U152 ( .A(n119), .B(n120), .C(n121), .Y(n31) );
  NAND2X1 U153 ( .A(n38), .B(n150), .Y(n121) );
  NAND3X1 U154 ( .A(n42), .B(n151), .C(n37), .Y(n150) );
  NAND2X1 U155 ( .A(B[7]), .B(A[7]), .Y(n37) );
  NAND3X1 U156 ( .A(n46), .B(n152), .C(n40), .Y(n151) );
  NAND2X1 U157 ( .A(n44), .B(n48), .Y(n152) );
  NAND2X1 U158 ( .A(B[4]), .B(A[4]), .Y(n48) );
  NAND2X1 U159 ( .A(B[5]), .B(A[5]), .Y(n44) );
  NAND2X1 U160 ( .A(B[6]), .B(A[6]), .Y(n42) );
  OR2X2 U161 ( .A(n153), .B(n154), .Y(n120) );
  NAND3X1 U162 ( .A(n46), .B(n49), .C(n40), .Y(n154) );
  OR2X2 U163 ( .A(A[6]), .B(B[6]), .Y(n40) );
  OR2X2 U164 ( .A(A[4]), .B(B[4]), .Y(n49) );
  OR2X2 U165 ( .A(A[5]), .B(B[5]), .Y(n46) );
  INVX2 U166 ( .A(n38), .Y(n153) );
  OR2X2 U167 ( .A(A[7]), .B(B[7]), .Y(n38) );
  INVX2 U168 ( .A(n155), .Y(n119) );
  OAI21X1 U169 ( .A(n156), .B(n157), .C(n54), .Y(n155) );
  NAND2X1 U170 ( .A(B[3]), .B(A[3]), .Y(n54) );
  OAI21X1 U171 ( .A(n158), .B(n159), .C(n53), .Y(n157) );
  OR2X2 U172 ( .A(A[3]), .B(B[3]), .Y(n53) );
  OAI21X1 U173 ( .A(n160), .B(n86), .C(n58), .Y(n159) );
  NAND2X1 U174 ( .A(B[2]), .B(A[2]), .Y(n58) );
  INVX2 U175 ( .A(n63), .Y(n160) );
  OR2X2 U176 ( .A(A[1]), .B(B[1]), .Y(n63) );
  INVX2 U177 ( .A(n61), .Y(n158) );
  NAND2X1 U178 ( .A(B[1]), .B(A[1]), .Y(n61) );
  INVX2 U179 ( .A(n56), .Y(n156) );
  OR2X2 U180 ( .A(A[2]), .B(B[2]), .Y(n56) );
  OR2X2 U181 ( .A(A[8]), .B(B[8]), .Y(n34) );
  NAND2X1 U182 ( .A(B[0]), .B(A[0]), .Y(n86) );
  OR2X2 U183 ( .A(A[0]), .B(B[0]), .Y(n87) );
endmodule


module matrix_math_DW01_add_12 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   \B[7] , \B[6] , \B[5] , \B[4] , \B[3] , \B[2] , \B[1] , \B[0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105;
  assign SUM[7] = \B[7] ;
  assign \B[7]  = B[7];
  assign SUM[6] = \B[6] ;
  assign \B[6]  = B[6];
  assign SUM[5] = \B[5] ;
  assign \B[5]  = B[5];
  assign SUM[4] = \B[4] ;
  assign \B[4]  = B[4];
  assign SUM[3] = \B[3] ;
  assign \B[3]  = B[3];
  assign SUM[2] = \B[2] ;
  assign \B[2]  = B[2];
  assign SUM[1] = \B[1] ;
  assign \B[1]  = B[1];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND2X1 U2 ( .A(n70), .B(n63), .Y(n69) );
  AND2X2 U3 ( .A(n94), .B(n95), .Y(n1) );
  NAND2X1 U4 ( .A(n30), .B(A[16]), .Y(n2) );
  OAI21X1 U5 ( .A(n41), .B(n42), .C(n43), .Y(n3) );
  INVX1 U6 ( .A(n53), .Y(n4) );
  INVX1 U7 ( .A(n53), .Y(n45) );
  OR2X2 U8 ( .A(n30), .B(A[16]), .Y(n70) );
  BUFX2 U9 ( .A(B[16]), .Y(n30) );
  OR2X2 U10 ( .A(B[20]), .B(A[20]), .Y(n5) );
  INVX1 U11 ( .A(n5), .Y(n6) );
  INVX1 U12 ( .A(n6), .Y(n7) );
  INVX1 U13 ( .A(n13), .Y(n8) );
  INVX2 U14 ( .A(n18), .Y(n13) );
  XOR2X1 U15 ( .A(n54), .B(n9), .Y(SUM[20]) );
  NAND2X1 U16 ( .A(n48), .B(n5), .Y(n9) );
  NOR2X1 U17 ( .A(B[22]), .B(A[22]), .Y(n10) );
  INVX1 U18 ( .A(n10), .Y(n39) );
  AND2X2 U19 ( .A(B[22]), .B(A[22]), .Y(n26) );
  BUFX4 U20 ( .A(B[16]), .Y(n31) );
  NAND2X1 U21 ( .A(n2), .B(n74), .Y(n11) );
  NAND2X1 U22 ( .A(n11), .B(n69), .Y(n68) );
  XOR2X1 U23 ( .A(n50), .B(n12), .Y(SUM[21]) );
  AND2X2 U24 ( .A(n44), .B(n43), .Y(n12) );
  INVX1 U25 ( .A(n8), .Y(n62) );
  INVX1 U26 ( .A(B[18]), .Y(n14) );
  INVX1 U27 ( .A(n14), .Y(n15) );
  INVX1 U28 ( .A(n17), .Y(n16) );
  AOI21X1 U29 ( .A(n58), .B(n57), .C(n59), .Y(n17) );
  NOR2X1 U30 ( .A(A[18]), .B(B[18]), .Y(n18) );
  INVX1 U31 ( .A(n96), .Y(n104) );
  AND2X1 U32 ( .A(n31), .B(A[16]), .Y(n28) );
  AND2X1 U33 ( .A(n32), .B(n35), .Y(SUM[8]) );
  XNOR2X1 U34 ( .A(n67), .B(n19), .Y(SUM[18]) );
  NAND2X1 U35 ( .A(n62), .B(n61), .Y(n19) );
  XNOR2X1 U36 ( .A(n45), .B(n56), .Y(SUM[19]) );
  XNOR2X1 U37 ( .A(n89), .B(n20), .Y(SUM[14]) );
  NAND2X1 U38 ( .A(n79), .B(n90), .Y(n20) );
  XOR2X1 U39 ( .A(n101), .B(n102), .Y(SUM[11]) );
  XOR2X1 U40 ( .A(n91), .B(n21), .Y(SUM[13]) );
  NAND2X1 U41 ( .A(n92), .B(n82), .Y(n21) );
  XNOR2X1 U42 ( .A(n1), .B(n22), .Y(SUM[12]) );
  NAND2X1 U43 ( .A(n84), .B(n85), .Y(n22) );
  XNOR2X1 U44 ( .A(n103), .B(n23), .Y(SUM[10]) );
  NAND2X1 U45 ( .A(n100), .B(n96), .Y(n23) );
  XOR2X1 U46 ( .A(n32), .B(n24), .Y(SUM[9]) );
  NAND2X1 U47 ( .A(n33), .B(n34), .Y(n24) );
  XOR2X1 U48 ( .A(n71), .B(n25), .Y(SUM[17]) );
  NAND2X1 U49 ( .A(n63), .B(n60), .Y(n25) );
  NOR2X1 U50 ( .A(A[15]), .B(B[15]), .Y(n27) );
  OR2X1 U51 ( .A(A[16]), .B(n31), .Y(n72) );
  XNOR2X1 U52 ( .A(n36), .B(n37), .Y(SUM[23]) );
  XOR2X1 U53 ( .A(B[23]), .B(A[23]), .Y(n37) );
  AOI21X1 U54 ( .A(n38), .B(n39), .C(n26), .Y(n36) );
  XOR2X1 U55 ( .A(n40), .B(n3), .Y(SUM[22]) );
  NOR2X1 U56 ( .A(n10), .B(n26), .Y(n40) );
  OAI21X1 U57 ( .A(n42), .B(n41), .C(n43), .Y(n38) );
  NAND2X1 U58 ( .A(n7), .B(n44), .Y(n42) );
  AOI21X1 U59 ( .A(n4), .B(n46), .C(n47), .Y(n41) );
  NAND2X1 U60 ( .A(n48), .B(n49), .Y(n47) );
  OR2X2 U61 ( .A(B[21]), .B(A[21]), .Y(n44) );
  NAND2X1 U62 ( .A(B[21]), .B(A[21]), .Y(n43) );
  NAND2X1 U63 ( .A(n48), .B(n51), .Y(n50) );
  NAND3X1 U64 ( .A(n46), .B(n5), .C(n52), .Y(n51) );
  NAND2X1 U65 ( .A(n53), .B(n49), .Y(n52) );
  NAND2X1 U66 ( .A(B[20]), .B(A[20]), .Y(n48) );
  AOI21X1 U67 ( .A(n16), .B(n46), .C(n55), .Y(n54) );
  INVX2 U68 ( .A(n49), .Y(n55) );
  NAND2X1 U69 ( .A(n49), .B(n46), .Y(n56) );
  OR2X2 U70 ( .A(A[19]), .B(B[19]), .Y(n46) );
  NAND2X1 U71 ( .A(B[19]), .B(A[19]), .Y(n49) );
  AOI21X1 U72 ( .A(n58), .B(n57), .C(n59), .Y(n53) );
  OAI21X1 U73 ( .A(n18), .B(n60), .C(n61), .Y(n59) );
  AND2X2 U74 ( .A(n13), .B(n63), .Y(n58) );
  AOI21X1 U75 ( .A(n64), .B(n74), .C(n65), .Y(n57) );
  NOR2X1 U76 ( .A(A[16]), .B(n31), .Y(n65) );
  NAND2X1 U77 ( .A(n31), .B(A[16]), .Y(n64) );
  NAND2X1 U78 ( .A(n15), .B(A[18]), .Y(n61) );
  NAND2X1 U79 ( .A(n60), .B(n68), .Y(n67) );
  NAND2X1 U80 ( .A(B[17]), .B(A[17]), .Y(n60) );
  OR2X2 U81 ( .A(B[17]), .B(A[17]), .Y(n63) );
  AOI21X1 U82 ( .A(n66), .B(n72), .C(n28), .Y(n71) );
  XNOR2X1 U83 ( .A(n73), .B(n74), .Y(SUM[16]) );
  INVX2 U84 ( .A(n66), .Y(n74) );
  OAI21X1 U85 ( .A(n27), .B(n75), .C(n76), .Y(n66) );
  OAI21X1 U86 ( .A(n77), .B(n78), .C(n79), .Y(n75) );
  OAI21X1 U87 ( .A(n80), .B(n81), .C(n82), .Y(n78) );
  OAI21X1 U88 ( .A(n83), .B(n1), .C(n84), .Y(n81) );
  INVX2 U89 ( .A(n85), .Y(n83) );
  XOR2X1 U90 ( .A(n31), .B(A[16]), .Y(n73) );
  XNOR2X1 U91 ( .A(n86), .B(n87), .Y(SUM[15]) );
  NOR2X1 U92 ( .A(n88), .B(n27), .Y(n87) );
  INVX2 U93 ( .A(n76), .Y(n88) );
  NAND2X1 U94 ( .A(B[15]), .B(A[15]), .Y(n76) );
  AOI21X1 U95 ( .A(n89), .B(n79), .C(n77), .Y(n86) );
  INVX2 U96 ( .A(n90), .Y(n77) );
  NAND2X1 U97 ( .A(B[14]), .B(A[14]), .Y(n90) );
  OR2X2 U98 ( .A(A[14]), .B(B[14]), .Y(n79) );
  OAI21X1 U99 ( .A(n80), .B(n91), .C(n82), .Y(n89) );
  INVX2 U100 ( .A(n92), .Y(n80) );
  NAND2X1 U101 ( .A(B[13]), .B(A[13]), .Y(n82) );
  OR2X2 U102 ( .A(A[13]), .B(B[13]), .Y(n92) );
  AND2X2 U103 ( .A(n93), .B(n85), .Y(n91) );
  NAND2X1 U104 ( .A(n1), .B(n84), .Y(n93) );
  NAND2X1 U105 ( .A(B[12]), .B(A[12]), .Y(n85) );
  OR2X2 U106 ( .A(A[12]), .B(B[12]), .Y(n84) );
  NAND3X1 U107 ( .A(n96), .B(n97), .C(n98), .Y(n95) );
  NAND3X1 U108 ( .A(n33), .B(n99), .C(n100), .Y(n97) );
  NAND2X1 U109 ( .A(n34), .B(n32), .Y(n99) );
  NAND2X1 U110 ( .A(n98), .B(n94), .Y(n102) );
  OR2X2 U111 ( .A(A[11]), .B(B[11]), .Y(n94) );
  NAND2X1 U112 ( .A(B[11]), .B(A[11]), .Y(n98) );
  AOI21X1 U113 ( .A(n103), .B(n100), .C(n104), .Y(n101) );
  NAND2X1 U114 ( .A(B[10]), .B(A[10]), .Y(n96) );
  OR2X2 U115 ( .A(A[10]), .B(B[10]), .Y(n100) );
  OAI21X1 U116 ( .A(n32), .B(n105), .C(n34), .Y(n103) );
  NAND2X1 U117 ( .A(B[9]), .B(A[9]), .Y(n34) );
  INVX2 U118 ( .A(n33), .Y(n105) );
  OR2X2 U119 ( .A(A[9]), .B(B[9]), .Y(n33) );
  NAND2X1 U120 ( .A(B[8]), .B(A[8]), .Y(n32) );
  OR2X2 U121 ( .A(A[8]), .B(B[8]), .Y(n35) );
endmodule


module matrix_math_DW01_add_18 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132;

  INVX1 U2 ( .A(A[19]), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(n22), .Y(n3) );
  BUFX2 U5 ( .A(n61), .Y(n4) );
  INVX1 U6 ( .A(n56), .Y(n13) );
  INVX1 U7 ( .A(n21), .Y(n5) );
  INVX2 U8 ( .A(A[18]), .Y(n21) );
  INVX1 U9 ( .A(n47), .Y(n6) );
  INVX1 U10 ( .A(n47), .Y(n33) );
  AND2X1 U11 ( .A(B[21]), .B(n8), .Y(n28) );
  INVX1 U12 ( .A(A[21]), .Y(n7) );
  INVX1 U13 ( .A(n7), .Y(n8) );
  OR2X2 U14 ( .A(A[19]), .B(B[19]), .Y(n9) );
  OR2X1 U15 ( .A(A[19]), .B(B[19]), .Y(n29) );
  AND2X1 U16 ( .A(B[19]), .B(A[19]), .Y(n64) );
  INVX1 U17 ( .A(A[20]), .Y(n10) );
  INVX1 U18 ( .A(A[20]), .Y(n23) );
  INVX1 U19 ( .A(n48), .Y(n11) );
  NAND2X1 U20 ( .A(n23), .B(n24), .Y(n12) );
  INVX2 U21 ( .A(B[20]), .Y(n24) );
  XOR2X1 U22 ( .A(n13), .B(n57), .Y(SUM[21]) );
  INVX2 U23 ( .A(n14), .Y(n44) );
  NAND3X1 U24 ( .A(n29), .B(n58), .C(n59), .Y(n14) );
  INVX2 U25 ( .A(n75), .Y(n19) );
  INVX2 U26 ( .A(n25), .Y(n26) );
  NAND2X1 U27 ( .A(B[7]), .B(A[7]), .Y(n15) );
  AND2X2 U28 ( .A(B[3]), .B(A[3]), .Y(n16) );
  NOR2X1 U29 ( .A(A[3]), .B(B[3]), .Y(n17) );
  NOR2X1 U30 ( .A(A[1]), .B(B[1]), .Y(n18) );
  XOR2X1 U31 ( .A(n76), .B(n19), .Y(SUM[18]) );
  XNOR2X1 U32 ( .A(n65), .B(n66), .Y(SUM[20]) );
  XOR2X1 U33 ( .A(n54), .B(n55), .Y(SUM[22]) );
  INVX1 U34 ( .A(n23), .Y(n20) );
  NAND2X1 U35 ( .A(n22), .B(n21), .Y(n73) );
  INVX1 U36 ( .A(B[18]), .Y(n22) );
  NAND2X1 U37 ( .A(n24), .B(n10), .Y(n58) );
  INVX1 U38 ( .A(B[20]), .Y(n25) );
  BUFX2 U39 ( .A(n62), .Y(n27) );
  AND2X1 U40 ( .A(B[17]), .B(A[17]), .Y(n74) );
  BUFX2 U41 ( .A(n5), .Y(n30) );
  BUFX2 U42 ( .A(n63), .Y(n31) );
  BUFX2 U43 ( .A(n3), .Y(n32) );
  XNOR2X1 U44 ( .A(n41), .B(n34), .Y(SUM[23]) );
  XNOR2X1 U45 ( .A(A[23]), .B(B[23]), .Y(n34) );
  INVX1 U46 ( .A(n48), .Y(n35) );
  NOR2X1 U47 ( .A(A[21]), .B(B[21]), .Y(n36) );
  INVX1 U48 ( .A(n36), .Y(n49) );
  AND2X1 U49 ( .A(n72), .B(n77), .Y(n37) );
  AND2X2 U50 ( .A(B[14]), .B(A[14]), .Y(n38) );
  AND2X2 U51 ( .A(B[12]), .B(A[12]), .Y(n39) );
  AND2X2 U52 ( .A(B[10]), .B(A[10]), .Y(n40) );
  AND2X1 U53 ( .A(n63), .B(n62), .Y(n60) );
  NAND2X1 U54 ( .A(n42), .B(n43), .Y(n41) );
  OAI21X1 U55 ( .A(n44), .B(n45), .C(n46), .Y(n43) );
  AOI21X1 U56 ( .A(n47), .B(n48), .C(n36), .Y(n46) );
  INVX2 U57 ( .A(B[22]), .Y(n48) );
  INVX2 U58 ( .A(A[22]), .Y(n47) );
  NAND3X1 U59 ( .A(n50), .B(n51), .C(n52), .Y(n45) );
  NAND2X1 U60 ( .A(A[21]), .B(B[21]), .Y(n51) );
  OAI21X1 U61 ( .A(n33), .B(n35), .C(n42), .Y(n55) );
  NAND2X1 U62 ( .A(n6), .B(n11), .Y(n42) );
  AOI21X1 U63 ( .A(n56), .B(n49), .C(n28), .Y(n54) );
  NAND2X1 U64 ( .A(n51), .B(n49), .Y(n57) );
  NAND3X1 U65 ( .A(n50), .B(n52), .C(n53), .Y(n56) );
  NAND3X1 U66 ( .A(n9), .B(n12), .C(n59), .Y(n53) );
  NAND2X1 U67 ( .A(n60), .B(n61), .Y(n59) );
  OAI21X1 U68 ( .A(A[20]), .B(B[20]), .C(n64), .Y(n50) );
  OAI21X1 U69 ( .A(n20), .B(n26), .C(n52), .Y(n66) );
  NAND2X1 U70 ( .A(A[20]), .B(B[20]), .Y(n52) );
  NAND2X1 U71 ( .A(n67), .B(n68), .Y(n65) );
  NAND2X1 U72 ( .A(n9), .B(n69), .Y(n68) );
  XNOR2X1 U73 ( .A(n70), .B(n69), .Y(SUM[19]) );
  NAND2X1 U74 ( .A(n67), .B(n9), .Y(n70) );
  NAND2X1 U75 ( .A(B[19]), .B(n2), .Y(n67) );
  NAND3X1 U76 ( .A(n31), .B(n27), .C(n4), .Y(n69) );
  NAND3X1 U77 ( .A(n71), .B(n72), .C(n73), .Y(n61) );
  OAI21X1 U78 ( .A(B[18]), .B(A[18]), .C(n74), .Y(n62) );
  OAI21X1 U79 ( .A(n30), .B(n32), .C(n31), .Y(n76) );
  NAND2X1 U80 ( .A(A[18]), .B(B[18]), .Y(n63) );
  NAND2X1 U81 ( .A(n77), .B(n78), .Y(n75) );
  NAND2X1 U82 ( .A(n71), .B(n72), .Y(n78) );
  NAND2X1 U83 ( .A(n79), .B(n80), .Y(n71) );
  OAI21X1 U84 ( .A(A[16]), .B(B[16]), .C(n81), .Y(n80) );
  NAND2X1 U85 ( .A(A[16]), .B(B[16]), .Y(n79) );
  XOR2X1 U86 ( .A(n82), .B(n37), .Y(SUM[17]) );
  NAND2X1 U87 ( .A(B[17]), .B(A[17]), .Y(n77) );
  OR2X2 U88 ( .A(B[17]), .B(A[17]), .Y(n72) );
  NAND2X1 U89 ( .A(n83), .B(n84), .Y(n82) );
  OAI21X1 U90 ( .A(B[16]), .B(A[16]), .C(n81), .Y(n84) );
  XNOR2X1 U91 ( .A(n81), .B(n85), .Y(SUM[16]) );
  OAI21X1 U92 ( .A(A[16]), .B(B[16]), .C(n83), .Y(n85) );
  NAND2X1 U93 ( .A(B[16]), .B(A[16]), .Y(n83) );
  OAI22X1 U94 ( .A(n86), .B(n87), .C(n88), .D(n89), .Y(n81) );
  OAI21X1 U95 ( .A(n38), .B(n90), .C(n91), .Y(n89) );
  OR2X2 U96 ( .A(A[14]), .B(B[14]), .Y(n91) );
  OAI21X1 U97 ( .A(n92), .B(n93), .C(n94), .Y(n90) );
  NAND2X1 U98 ( .A(B[13]), .B(A[13]), .Y(n94) );
  OAI21X1 U99 ( .A(n39), .B(n95), .C(n96), .Y(n93) );
  OR2X2 U100 ( .A(A[12]), .B(B[12]), .Y(n96) );
  OAI22X1 U101 ( .A(n97), .B(n98), .C(n99), .D(n100), .Y(n95) );
  OAI21X1 U102 ( .A(n101), .B(n40), .C(n102), .Y(n100) );
  OR2X2 U103 ( .A(A[10]), .B(B[10]), .Y(n102) );
  NAND3X1 U104 ( .A(n103), .B(n104), .C(n105), .Y(n101) );
  NAND2X1 U105 ( .A(B[9]), .B(A[9]), .Y(n105) );
  NAND3X1 U106 ( .A(n106), .B(n107), .C(n108), .Y(n104) );
  AOI22X1 U107 ( .A(n109), .B(n110), .C(n111), .D(n112), .Y(n107) );
  INVX2 U108 ( .A(A[8]), .Y(n112) );
  INVX2 U109 ( .A(B[8]), .Y(n111) );
  INVX2 U110 ( .A(A[7]), .Y(n110) );
  INVX2 U111 ( .A(B[7]), .Y(n109) );
  NAND3X1 U112 ( .A(n113), .B(n114), .C(n15), .Y(n106) );
  OAI21X1 U113 ( .A(n117), .B(n16), .C(n115), .Y(n114) );
  INVX2 U114 ( .A(n118), .Y(n115) );
  NAND3X1 U115 ( .A(n119), .B(n120), .C(n121), .Y(n118) );
  OR2X2 U116 ( .A(A[4]), .B(B[4]), .Y(n119) );
  AOI21X1 U117 ( .A(n122), .B(n123), .C(n17), .Y(n117) );
  NAND2X1 U118 ( .A(n124), .B(n116), .Y(n123) );
  OR2X2 U119 ( .A(A[2]), .B(B[2]), .Y(n116) );
  OAI22X1 U120 ( .A(n125), .B(n126), .C(n18), .D(n127), .Y(n124) );
  NAND2X1 U121 ( .A(A[0]), .B(B[0]), .Y(n127) );
  INVX2 U122 ( .A(B[1]), .Y(n126) );
  INVX2 U123 ( .A(A[1]), .Y(n125) );
  NAND2X1 U124 ( .A(B[2]), .B(A[2]), .Y(n122) );
  AOI22X1 U125 ( .A(B[6]), .B(A[6]), .C(n128), .D(n121), .Y(n113) );
  OR2X2 U126 ( .A(A[6]), .B(B[6]), .Y(n121) );
  AOI21X1 U127 ( .A(n129), .B(n130), .C(n131), .Y(n128) );
  INVX2 U128 ( .A(n120), .Y(n131) );
  OR2X2 U129 ( .A(A[5]), .B(B[5]), .Y(n120) );
  NAND2X1 U130 ( .A(B[5]), .B(A[5]), .Y(n130) );
  NAND2X1 U131 ( .A(B[4]), .B(A[4]), .Y(n129) );
  NAND2X1 U132 ( .A(n132), .B(n108), .Y(n103) );
  OR2X2 U133 ( .A(A[9]), .B(B[9]), .Y(n108) );
  AND2X2 U134 ( .A(A[8]), .B(B[8]), .Y(n132) );
  NOR2X1 U135 ( .A(A[11]), .B(B[11]), .Y(n99) );
  INVX2 U136 ( .A(B[11]), .Y(n98) );
  INVX2 U137 ( .A(A[11]), .Y(n97) );
  NOR2X1 U138 ( .A(A[13]), .B(B[13]), .Y(n92) );
  NOR2X1 U139 ( .A(A[15]), .B(B[15]), .Y(n88) );
  INVX2 U140 ( .A(B[15]), .Y(n87) );
  INVX2 U141 ( .A(A[15]), .Y(n86) );
endmodule


module matrix_math ( screen_cor, init_matrix, clk, rst_n, row_sel, sel, 
        math_done, strb_screen, point, row, err );
  output [7:0] screen_cor;
  output [1:0] row_sel;
  input [47:0] point;
  input [63:0] row;
  input init_matrix, clk, rst_n;
  output sel, math_done, strb_screen, err;
  wire   \V1[23] , n32, n33, n34, n35, N99, N98, N97, N96, N95, N94, N93, N92,
         N91, N90, N9, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N8,
         N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N7, N69, N68, N67,
         N66, N65, N64, N63, N62, N61, N60, N6, N59, N58, N57, N56, N55, N54,
         N53, N52, N51, N50, N5, N49, N48, N47, N46, N45, N44, N43, N42, N41,
         N40, N4, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N3, N29,
         N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19, N18, N17, N16,
         N15, N14, N13, N12, N119, N118, N117, N116, N115, N114, N113, N112,
         N111, N110, N11, N109, N108, N107, N106, N105, N104, N103, N102, N101,
         N100, N10, N1, N0, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n48;
  wire   [3:0] state;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39;
  assign err = 1'b0;
  assign row_sel[1] = 1'b0;

  DFFSR \state_reg[0]  ( .D(n48), .CLK(clk), .R(rst_n), .S(1'b1), .Q(state[0])
         );
  DFFSR \state_reg[1]  ( .D(n34), .CLK(clk), .R(rst_n), .S(1'b1), .Q(state[1])
         );
  DFFSR \state_reg[2]  ( .D(n33), .CLK(clk), .R(rst_n), .S(1'b1), .Q(state[2])
         );
  DFFSR \state_reg[3]  ( .D(n14), .CLK(clk), .R(rst_n), .S(1'b1), .Q(state[3])
         );
  NAND2X1 U39 ( .A(n18), .B(n12), .Y(n32) );
  matrix_math_DW02_mult_2 mult_53 ( .A(row[63:48]), .B(point[47:32]), .TC(1'b1), .PRODUCT({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
        N4, N3, N2, N1, N0}) );
  matrix_math_DW02_mult_1 mult_53_2 ( .A(row[47:32]), .B(point[31:16]), .TC(
        1'b1), .PRODUCT({SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24}) );
  matrix_math_DW02_mult_0 mult_53_3 ( .A(row[31:16]), .B(point[15:0]), .TC(
        1'b1), .PRODUCT({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, N95, N94, N93, N92, 
        N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, 
        N77, N76, N75, N74, N73, N72}) );
  matrix_math_DW01_add_13 add_1_root_add_0_root_add_53_3 ( .A({N23, N22, N21, 
        N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, 
        N5, N4, N3, N2, N1, N0}), .B({N95, N94, N93, N92, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, 
        N73, N72}), .CI(1'b0), .SUM({N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48}) );
  matrix_math_DW01_add_12 add_2_root_add_0_root_add_53_3 ( .A({row[15:0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24}), .CI(1'b0), .SUM({N119, N118, N117, 
        N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, 
        N104, N103, N102, N101, N100, N99, N98, N97, N96}) );
  matrix_math_DW01_add_18 add_0_root_add_0_root_add_53_3 ( .A({N71, N70, N69, 
        N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50, N49, N48}), .B({N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96}), .CI(1'b0), .SUM({\V1[23] , 
        screen_cor[6:0], SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39}) );
  BUFX2 U6 ( .A(n22), .Y(n5) );
  BUFX2 U7 ( .A(state[1]), .Y(n6) );
  INVX1 U8 ( .A(state[1]), .Y(n17) );
  BUFX4 U9 ( .A(state[0]), .Y(n7) );
  BUFX2 U10 ( .A(state[0]), .Y(n16) );
  INVX2 U11 ( .A(n17), .Y(n8) );
  INVX1 U12 ( .A(n28), .Y(n9) );
  INVX1 U13 ( .A(n35), .Y(n36) );
  INVX2 U14 ( .A(state[2]), .Y(n10) );
  INVX4 U15 ( .A(n10), .Y(n11) );
  BUFX4 U16 ( .A(state[3]), .Y(n12) );
  INVX1 U17 ( .A(state[3]), .Y(n39) );
  BUFX2 U18 ( .A(n8), .Y(n13) );
  OAI21X1 U19 ( .A(n24), .B(n23), .C(n22), .Y(n14) );
  INVX2 U20 ( .A(n15), .Y(strb_screen) );
  AND2X2 U21 ( .A(n21), .B(n5), .Y(n15) );
  BUFX2 U22 ( .A(n7), .Y(n18) );
  INVX1 U23 ( .A(n6), .Y(n24) );
  OR2X2 U24 ( .A(n18), .B(n12), .Y(n46) );
  INVX2 U25 ( .A(n46), .Y(n41) );
  OR2X2 U26 ( .A(n13), .B(n11), .Y(n38) );
  NAND2X1 U27 ( .A(n41), .B(n38), .Y(n21) );
  INVX2 U28 ( .A(n11), .Y(n29) );
  NOR2X1 U29 ( .A(n6), .B(n16), .Y(n20) );
  NAND3X1 U30 ( .A(n12), .B(n29), .C(n20), .Y(n22) );
  NOR2X1 U31 ( .A(n32), .B(n38), .Y(math_done) );
  NAND3X1 U32 ( .A(n11), .B(n7), .C(n39), .Y(n23) );
  OAI21X1 U33 ( .A(n24), .B(n23), .C(n22), .Y(n35) );
  NAND2X1 U34 ( .A(n6), .B(n16), .Y(n25) );
  NOR2X1 U35 ( .A(n12), .B(n25), .Y(n27) );
  NOR3X1 U36 ( .A(n7), .B(n12), .C(n8), .Y(n26) );
  MUX2X1 U37 ( .B(n27), .A(n26), .S(n11), .Y(n37) );
  INVX2 U38 ( .A(n37), .Y(n28) );
  OR2X2 U40 ( .A(n28), .B(n14), .Y(sel) );
  NOR2X1 U41 ( .A(n12), .B(n29), .Y(n31) );
  XOR2X1 U42 ( .A(n7), .B(n8), .Y(n30) );
  NAND2X1 U43 ( .A(n31), .B(n30), .Y(n43) );
  NAND2X1 U44 ( .A(n36), .B(n43), .Y(row_sel[0]) );
  INVX2 U45 ( .A(\V1[23] ), .Y(screen_cor[7]) );
  NAND2X1 U46 ( .A(n43), .B(n9), .Y(n33) );
  INVX2 U47 ( .A(n38), .Y(n40) );
  NAND3X1 U48 ( .A(n18), .B(n40), .C(n39), .Y(n44) );
  NAND2X1 U49 ( .A(n13), .B(n41), .Y(n42) );
  NAND3X1 U50 ( .A(n44), .B(n43), .C(n42), .Y(n34) );
  INVX2 U51 ( .A(init_matrix), .Y(n45) );
  OAI21X1 U52 ( .A(n46), .B(n45), .C(n15), .Y(n48) );
endmodule


module Rasterizer_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module Rasterizer_DW01_add_0 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [11:1] carry;

  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X2 U2 ( .A(carry[9]), .B(A[9]), .Y(n2) );
  AND2X2 U3 ( .A(n2), .B(A[10]), .Y(n3) );
  XOR2X1 U4 ( .A(A[11]), .B(n3), .Y(SUM[11]) );
  XOR2X1 U5 ( .A(n2), .B(A[10]), .Y(SUM[10]) );
  XOR2X1 U6 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  XOR2X1 U7 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Rasterizer_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module Rasterizer_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [12:0] carry;

  FAX1 U2_8 ( .A(A[8]), .B(n9), .C(carry[8]), .YC(carry[9]), .YS(DIFF[8]) );
  FAX1 U2_7 ( .A(A[7]), .B(n8), .C(carry[7]), .YC(carry[8]), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n7), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n6), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n5), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n4), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n3), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n2), .C(carry[1]), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X2 U1 ( .A(A[10]), .B(carry[10]), .Y(carry[11]) );
  XNOR2X1 U2 ( .A(carry[10]), .B(A[10]), .Y(DIFF[10]) );
  XNOR2X1 U3 ( .A(A[11]), .B(carry[11]), .Y(DIFF[11]) );
  OR2X2 U4 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
  XNOR2X1 U5 ( .A(carry[9]), .B(A[9]), .Y(DIFF[9]) );
  OR2X2 U6 ( .A(A[0]), .B(n1), .Y(carry[1]) );
  XNOR2X1 U7 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
  INVX2 U8 ( .A(B[0]), .Y(n1) );
  INVX2 U9 ( .A(B[1]), .Y(n2) );
  INVX2 U10 ( .A(B[2]), .Y(n3) );
  INVX2 U11 ( .A(B[3]), .Y(n4) );
  INVX2 U12 ( .A(B[4]), .Y(n5) );
  INVX2 U13 ( .A(B[5]), .Y(n6) );
  INVX2 U14 ( .A(B[6]), .Y(n7) );
  INVX2 U15 ( .A(B[7]), .Y(n8) );
  INVX2 U16 ( .A(B[8]), .Y(n9) );
endmodule


module Rasterizer_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module Rasterizer_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n1), .C(carry[7]), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n2), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n3), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n4), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n5), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n6), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n7), .C(carry[1]), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X2 U1 ( .A(A[0]), .B(n8), .Y(carry[1]) );
  XNOR2X1 U2 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  INVX2 U3 ( .A(B[7]), .Y(n1) );
  INVX2 U4 ( .A(B[6]), .Y(n2) );
  INVX2 U5 ( .A(B[5]), .Y(n3) );
  INVX2 U6 ( .A(B[4]), .Y(n4) );
  INVX2 U7 ( .A(B[3]), .Y(n5) );
  INVX2 U8 ( .A(B[2]), .Y(n6) );
  INVX2 U9 ( .A(B[1]), .Y(n7) );
  INVX2 U10 ( .A(B[0]), .Y(n8) );
endmodule


module Rasterizer_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n1), .C(carry[7]), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n2), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n3), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n4), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n5), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n6), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n7), .C(carry[1]), .YC(carry[2]), .YS(DIFF[1]) );
  INVX1 U1 ( .A(B[7]), .Y(n1) );
  OR2X2 U2 ( .A(A[0]), .B(n8), .Y(carry[1]) );
  XNOR2X1 U3 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  INVX2 U4 ( .A(B[6]), .Y(n2) );
  INVX2 U5 ( .A(B[5]), .Y(n3) );
  INVX2 U6 ( .A(B[4]), .Y(n4) );
  INVX2 U7 ( .A(B[3]), .Y(n5) );
  INVX2 U8 ( .A(B[2]), .Y(n6) );
  INVX2 U9 ( .A(B[1]), .Y(n7) );
  INVX2 U10 ( .A(B[0]), .Y(n8) );
endmodule


module Rasterizer_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n1), .C(carry[7]), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n2), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n3), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n4), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n5), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n6), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n7), .C(carry[1]), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X2 U1 ( .A(A[0]), .B(n8), .Y(carry[1]) );
  XNOR2X1 U2 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  INVX2 U3 ( .A(B[7]), .Y(n1) );
  INVX2 U4 ( .A(B[6]), .Y(n2) );
  INVX2 U5 ( .A(B[5]), .Y(n3) );
  INVX2 U6 ( .A(B[4]), .Y(n4) );
  INVX2 U7 ( .A(B[3]), .Y(n5) );
  INVX2 U8 ( .A(B[2]), .Y(n6) );
  INVX2 U9 ( .A(B[1]), .Y(n7) );
  INVX2 U10 ( .A(B[0]), .Y(n8) );
endmodule


module Rasterizer_DW01_sub_6 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n1), .C(carry[7]), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n2), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n3), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n4), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n5), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n6), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n7), .C(carry[1]), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X2 U1 ( .A(A[0]), .B(n8), .Y(carry[1]) );
  XNOR2X1 U2 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  INVX2 U3 ( .A(B[7]), .Y(n1) );
  INVX2 U4 ( .A(B[6]), .Y(n2) );
  INVX2 U5 ( .A(B[5]), .Y(n3) );
  INVX2 U6 ( .A(B[4]), .Y(n4) );
  INVX2 U7 ( .A(B[3]), .Y(n5) );
  INVX2 U8 ( .A(B[2]), .Y(n6) );
  INVX2 U9 ( .A(B[1]), .Y(n7) );
  INVX2 U10 ( .A(B[0]), .Y(n8) );
endmodule


module Rasterizer_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [8:1] carry;

  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Rasterizer ( clk, X0, X1, Y0, Y1, init_rast, RST_N, rast_done, 
        rast_strb, rast_index, rast_addr );
  input [7:0] X0;
  input [7:0] X1;
  input [7:0] Y0;
  input [7:0] Y1;
  output [3:0] rast_index;
  output [15:0] rast_addr;
  input clk, init_rast, RST_N;
  output rast_done, rast_strb;
  wire   iX, iY, steep, N95, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N121, N123, N124, N125,
         N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N188, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, N229, N230, N231, N232, N257, N258, N259, N260, N261,
         N262, N263, N264, N265, N266, N269, N270, N271, N272, N273, N274,
         N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285,
         N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296,
         N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316,
         N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327,
         N328, N329, N330, N331, N332, N333, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, N198, N197, N196,
         N195, N194, N193, N192, N191, N190,
         \sub_1_root_sub_0_root_sub_184/carry[7] ,
         \sub_1_root_sub_0_root_sub_184/carry[6] ,
         \sub_1_root_sub_0_root_sub_184/carry[5] ,
         \sub_1_root_sub_0_root_sub_184/carry[4] ,
         \sub_1_root_sub_0_root_sub_184/carry[3] ,
         \sub_1_root_sub_0_root_sub_184/carry[2] , n1, n2, n5, n6, n7, n8, n9,
         n10, n11, n12, n15, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n264, n265, n361, n362, n398, n399, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642;
  wire   [3:0] state;
  wire   [8:0] dx;
  wire   [8:0] dy;
  wire   [11:0] err;
  wire   [7:0] i;
  wire   [3:0] count;
  wire   [3:0] nextstate;
  assign rast_addr[12] = 1'b0;
  assign rast_addr[13] = 1'b0;
  assign rast_addr[14] = 1'b0;
  assign rast_addr[15] = 1'b0;

  DFFSR \i_reg[0]  ( .D(n567), .CLK(clk), .R(n24), .S(1'b1), .Q(i[0]) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n21), .S(1'b1), .Q(
        state[2]) );
  DFFSR \dx_reg[0]  ( .D(n529), .CLK(clk), .R(n21), .S(1'b1), .Q(dx[0]) );
  DFFSR \dx_reg[1]  ( .D(n528), .CLK(clk), .R(n21), .S(1'b1), .Q(N190) );
  DFFSR \dx_reg[2]  ( .D(n527), .CLK(clk), .R(n21), .S(1'b1), .Q(dx[2]) );
  DFFSR \dx_reg[3]  ( .D(n526), .CLK(clk), .R(n21), .S(1'b1), .Q(dx[3]) );
  DFFSR \dx_reg[4]  ( .D(n525), .CLK(clk), .R(n21), .S(1'b1), .Q(dx[4]) );
  DFFSR \dx_reg[5]  ( .D(n524), .CLK(clk), .R(n21), .S(1'b1), .Q(dx[5]) );
  DFFSR \dx_reg[6]  ( .D(n523), .CLK(clk), .R(n21), .S(1'b1), .Q(dx[6]) );
  DFFSR \dx_reg[7]  ( .D(n522), .CLK(clk), .R(n21), .S(1'b1), .Q(dx[7]) );
  DFFSR \dx_reg[8]  ( .D(n521), .CLK(clk), .R(n21), .S(1'b1), .Q(dx[8]) );
  DFFSR \dy_reg[8]  ( .D(n530), .CLK(clk), .R(n21), .S(1'b1), .Q(dy[8]) );
  DFFSR \dy_reg[7]  ( .D(n531), .CLK(clk), .R(n22), .S(1'b1), .Q(dy[7]) );
  DFFSR \err_reg[11]  ( .D(n554), .CLK(clk), .R(n22), .S(1'b1), .Q(err[11]) );
  DFFSR \err_reg[10]  ( .D(n549), .CLK(clk), .R(n22), .S(1'b1), .Q(err[10]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n22), .S(1'b1), .Q(
        state[1]) );
  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n22), .S(1'b1), .Q(
        state[0]) );
  DFFSR \count_reg[3]  ( .D(n550), .CLK(clk), .R(n22), .S(1'b1), .Q(count[3])
         );
  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(clk), .R(n22), .S(1'b1), .Q(
        state[3]) );
  DFFSR \dy_reg[0]  ( .D(n538), .CLK(clk), .R(n22), .S(1'b1), .Q(dy[0]) );
  DFFSR \dy_reg[1]  ( .D(n537), .CLK(clk), .R(n22), .S(1'b1), .Q(dy[1]) );
  DFFSR \dy_reg[2]  ( .D(n536), .CLK(clk), .R(n22), .S(1'b1), .Q(dy[2]) );
  DFFSR \dy_reg[3]  ( .D(n535), .CLK(clk), .R(n22), .S(1'b1), .Q(dy[3]) );
  DFFSR \dy_reg[4]  ( .D(n534), .CLK(clk), .R(n22), .S(1'b1), .Q(dy[4]) );
  DFFSR \dy_reg[5]  ( .D(n533), .CLK(clk), .R(n23), .S(1'b1), .Q(dy[5]) );
  DFFSR \dy_reg[6]  ( .D(n532), .CLK(clk), .R(n23), .S(1'b1), .Q(dy[6]) );
  DFFSR \count_reg[0]  ( .D(n553), .CLK(clk), .R(n23), .S(1'b1), .Q(count[0])
         );
  DFFSR \count_reg[1]  ( .D(n552), .CLK(clk), .R(n23), .S(1'b1), .Q(count[1])
         );
  DFFSR \count_reg[2]  ( .D(n551), .CLK(clk), .R(n23), .S(1'b1), .Q(count[2])
         );
  DFFSR iX_reg ( .D(n519), .CLK(clk), .R(n23), .S(1'b1), .Q(iX) );
  DFFSR iY_reg ( .D(n520), .CLK(clk), .R(n23), .S(1'b1), .Q(iY) );
  DFFSR \err_reg[9]  ( .D(n548), .CLK(clk), .R(n23), .S(1'b1), .Q(err[9]) );
  DFFSR \err_reg[8]  ( .D(n555), .CLK(clk), .R(1'b1), .S(n27), .Q(err[8]) );
  DFFSR \err_reg[7]  ( .D(n547), .CLK(clk), .R(n23), .S(1'b1), .Q(err[7]) );
  DFFSR \err_reg[6]  ( .D(n546), .CLK(clk), .R(n23), .S(1'b1), .Q(err[6]) );
  DFFSR \err_reg[5]  ( .D(n545), .CLK(clk), .R(n23), .S(1'b1), .Q(err[5]) );
  DFFSR \err_reg[4]  ( .D(n544), .CLK(clk), .R(n23), .S(1'b1), .Q(err[4]) );
  DFFSR \err_reg[3]  ( .D(n543), .CLK(clk), .R(n24), .S(1'b1), .Q(err[3]) );
  DFFSR \err_reg[2]  ( .D(n542), .CLK(clk), .R(n24), .S(1'b1), .Q(err[2]) );
  DFFSR \err_reg[1]  ( .D(n541), .CLK(clk), .R(n24), .S(1'b1), .Q(err[1]) );
  DFFSR \err_reg[0]  ( .D(n540), .CLK(clk), .R(n24), .S(1'b1), .Q(err[0]) );
  DFFSR steep_reg ( .D(n539), .CLK(clk), .R(n24), .S(1'b1), .Q(steep) );
  DFFSR \Y_reg[0]  ( .D(n518), .CLK(clk), .R(n24), .S(1'b1), .Q(N213) );
  DFFSR \X_reg[0]  ( .D(n510), .CLK(clk), .R(n24), .S(1'b1), .Q(N229) );
  DFFSR \X_reg[7]  ( .D(n499), .CLK(clk), .R(n24), .S(1'b1), .Q(N212) );
  DFFSR \Y_reg[7]  ( .D(n511), .CLK(clk), .R(n24), .S(1'b1), .Q(N220) );
  DFFSR \Y_reg[6]  ( .D(n512), .CLK(clk), .R(n24), .S(1'b1), .Q(N219) );
  DFFSR \X_reg[6]  ( .D(n500), .CLK(clk), .R(n24), .S(1'b1), .Q(N211) );
  DFFSR \X_reg[5]  ( .D(n501), .CLK(clk), .R(n25), .S(1'b1), .Q(N210) );
  DFFSR \Y_reg[5]  ( .D(n513), .CLK(clk), .R(n25), .S(1'b1), .Q(N218) );
  DFFSR \Y_reg[1]  ( .D(n517), .CLK(clk), .R(n25), .S(1'b1), .Q(N214) );
  DFFSR \X_reg[1]  ( .D(n509), .CLK(clk), .R(n25), .S(1'b1), .Q(N230) );
  DFFSR \rast_indexi_reg[1]  ( .D(n505), .CLK(clk), .R(n25), .S(1'b1), .Q(
        rast_index[1]) );
  DFFSR \Y_reg[2]  ( .D(n516), .CLK(clk), .R(n25), .S(1'b1), .Q(N215) );
  DFFSR \X_reg[2]  ( .D(n508), .CLK(clk), .R(n25), .S(1'b1), .Q(N231) );
  DFFSR \rast_indexi_reg[2]  ( .D(n504), .CLK(clk), .R(n25), .S(1'b1), .Q(
        rast_index[2]) );
  DFFSR \Y_reg[3]  ( .D(n515), .CLK(clk), .R(n25), .S(1'b1), .Q(N216) );
  DFFSR \X_reg[3]  ( .D(n507), .CLK(clk), .R(n25), .S(1'b1), .Q(N232) );
  DFFSR \rast_indexi_reg[3]  ( .D(n503), .CLK(clk), .R(n25), .S(1'b1), .Q(
        rast_index[3]) );
  DFFSR \Y_reg[4]  ( .D(n514), .CLK(clk), .R(n26), .S(1'b1), .Q(N217) );
  DFFSR \X_reg[4]  ( .D(n502), .CLK(clk), .R(n26), .S(1'b1), .Q(N209) );
  DFFSR \rast_addri_reg[4]  ( .D(n498), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[0]) );
  DFFSR \rast_addri_reg[5]  ( .D(n497), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[1]) );
  DFFSR \rast_addri_reg[6]  ( .D(n496), .CLK(clk), .R(n25), .S(1'b1), .Q(
        rast_addr[2]) );
  DFFSR \rast_addri_reg[7]  ( .D(n495), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[3]) );
  DFFSR \rast_addri_reg[8]  ( .D(n494), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[4]) );
  DFFSR \rast_addri_reg[9]  ( .D(n493), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[5]) );
  DFFSR \rast_addri_reg[10]  ( .D(n492), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[6]) );
  DFFSR \rast_addri_reg[11]  ( .D(n491), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[7]) );
  DFFSR \rast_addri_reg[12]  ( .D(n490), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[8]) );
  DFFSR \rast_addri_reg[13]  ( .D(n489), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[9]) );
  DFFSR \rast_addri_reg[14]  ( .D(n488), .CLK(clk), .R(n26), .S(1'b1), .Q(
        rast_addr[10]) );
  DFFSR \rast_addri_reg[15]  ( .D(n487), .CLK(clk), .R(n27), .S(1'b1), .Q(
        rast_addr[11]) );
  DFFSR \rast_indexi_reg[0]  ( .D(n506), .CLK(clk), .R(n27), .S(1'b1), .Q(
        rast_index[0]) );
  DFFSR \i_reg[7]  ( .D(n568), .CLK(clk), .R(n27), .S(1'b1), .Q(i[7]) );
  DFFSR \i_reg[1]  ( .D(n574), .CLK(clk), .R(n27), .S(1'b1), .Q(i[1]) );
  DFFSR \i_reg[2]  ( .D(n573), .CLK(clk), .R(n27), .S(1'b1), .Q(i[2]) );
  DFFSR \i_reg[3]  ( .D(n572), .CLK(clk), .R(n27), .S(1'b1), .Q(i[3]) );
  DFFSR \i_reg[4]  ( .D(n571), .CLK(clk), .R(n27), .S(1'b1), .Q(i[4]) );
  DFFSR \i_reg[5]  ( .D(n570), .CLK(clk), .R(n27), .S(1'b1), .Q(i[5]) );
  DFFSR \i_reg[6]  ( .D(n569), .CLK(clk), .R(n21), .S(1'b1), .Q(i[6]) );
  AND2X2 U102 ( .A(n255), .B(n256), .Y(n249) );
  OR2X2 U104 ( .A(n312), .B(n612), .Y(n281) );
  OR2X2 U105 ( .A(n312), .B(n611), .Y(n317) );
  AND2X2 U106 ( .A(state[1]), .B(n616), .Y(n477) );
  AND2X2 U107 ( .A(state[1]), .B(state[0]), .Y(n484) );
  NOR2X1 U188 ( .A(n229), .B(n230), .Y(rast_strb) );
  NAND2X1 U189 ( .A(n599), .B(n621), .Y(n230) );
  NAND3X1 U190 ( .A(n623), .B(n618), .C(n622), .Y(n229) );
  NAND3X1 U191 ( .A(n598), .B(n231), .C(n232), .Y(nextstate[3]) );
  NOR2X1 U192 ( .A(n612), .B(n233), .Y(n232) );
  NAND2X1 U193 ( .A(n234), .B(n235), .Y(n233) );
  OAI21X1 U194 ( .A(count[2]), .B(n236), .C(n599), .Y(n231) );
  NAND3X1 U195 ( .A(n237), .B(n598), .C(n238), .Y(nextstate[2]) );
  NOR2X1 U196 ( .A(n239), .B(n240), .Y(n238) );
  NAND2X1 U197 ( .A(n241), .B(n242), .Y(n240) );
  NAND2X1 U198 ( .A(n243), .B(n244), .Y(n239) );
  OAI21X1 U199 ( .A(n246), .B(n247), .C(n248), .Y(n245) );
  NOR2X1 U200 ( .A(n236), .B(n623), .Y(n246) );
  AOI21X1 U201 ( .A(N265), .B(n601), .C(n611), .Y(n237) );
  NAND3X1 U202 ( .A(n249), .B(n250), .C(n251), .Y(nextstate[1]) );
  NOR2X1 U203 ( .A(n610), .B(n252), .Y(n251) );
  OAI21X1 U204 ( .A(N266), .B(n234), .C(n253), .Y(n252) );
  NAND3X1 U205 ( .A(n599), .B(n623), .C(n617), .Y(n253) );
  NAND3X1 U206 ( .A(n622), .B(n618), .C(count[0]), .Y(n236) );
  NOR2X1 U207 ( .A(n603), .B(n606), .Y(n250) );
  NAND3X1 U208 ( .A(n257), .B(n258), .C(n259), .Y(nextstate[0]) );
  NOR2X1 U209 ( .A(n260), .B(n261), .Y(n259) );
  NAND2X1 U210 ( .A(n262), .B(n243), .Y(n261) );
  NAND2X1 U211 ( .A(n248), .B(n244), .Y(n260) );
  AOI21X1 U212 ( .A(init_rast), .B(n608), .C(n605), .Y(n258) );
  AOI22X1 U213 ( .A(N266), .B(n609), .C(n607), .D(n613), .Y(n257) );
  OAI21X1 U214 ( .A(n576), .B(n641), .C(n263), .Y(n487) );
  AOI22X1 U215 ( .A(N220), .B(n9), .C(N212), .D(n1), .Y(n263) );
  OAI21X1 U216 ( .A(n576), .B(n640), .C(n266), .Y(n488) );
  AOI22X1 U217 ( .A(N219), .B(n9), .C(N211), .D(n1), .Y(n266) );
  OAI21X1 U218 ( .A(n576), .B(n639), .C(n267), .Y(n489) );
  AOI22X1 U219 ( .A(N218), .B(n9), .C(N210), .D(n1), .Y(n267) );
  OAI21X1 U220 ( .A(n576), .B(n638), .C(n268), .Y(n490) );
  AOI22X1 U221 ( .A(N217), .B(n9), .C(N209), .D(n1), .Y(n268) );
  OAI21X1 U222 ( .A(n576), .B(n637), .C(n269), .Y(n491) );
  AOI22X1 U223 ( .A(N216), .B(n9), .C(N232), .D(n1), .Y(n269) );
  OAI21X1 U224 ( .A(n576), .B(n636), .C(n270), .Y(n492) );
  AOI22X1 U225 ( .A(N215), .B(n9), .C(N231), .D(n1), .Y(n270) );
  OAI21X1 U226 ( .A(n576), .B(n635), .C(n271), .Y(n493) );
  AOI22X1 U227 ( .A(N214), .B(n9), .C(N230), .D(n1), .Y(n271) );
  OAI21X1 U228 ( .A(n576), .B(n634), .C(n272), .Y(n494) );
  AOI22X1 U229 ( .A(N213), .B(n9), .C(N229), .D(n1), .Y(n272) );
  OAI21X1 U230 ( .A(n576), .B(n633), .C(n273), .Y(n495) );
  AOI22X1 U231 ( .A(N212), .B(n9), .C(N220), .D(n1), .Y(n273) );
  OAI21X1 U232 ( .A(n576), .B(n632), .C(n274), .Y(n496) );
  AOI22X1 U233 ( .A(N211), .B(n9), .C(N219), .D(n1), .Y(n274) );
  OAI21X1 U234 ( .A(n576), .B(n631), .C(n275), .Y(n497) );
  AOI22X1 U235 ( .A(N210), .B(n9), .C(N218), .D(n1), .Y(n275) );
  OAI21X1 U236 ( .A(n576), .B(n630), .C(n276), .Y(n498) );
  AOI22X1 U237 ( .A(N209), .B(n9), .C(N217), .D(n1), .Y(n276) );
  NAND3X1 U238 ( .A(n277), .B(n278), .C(n279), .Y(n499) );
  AOI22X1 U239 ( .A(N333), .B(n280), .C(N212), .D(n281), .Y(n279) );
  NAND2X1 U240 ( .A(N325), .B(n282), .Y(n278) );
  AOI22X1 U241 ( .A(N220), .B(n283), .C(X0[7]), .D(n606), .Y(n277) );
  NAND3X1 U242 ( .A(n284), .B(n285), .C(n286), .Y(n500) );
  AOI22X1 U243 ( .A(N332), .B(n280), .C(N211), .D(n281), .Y(n286) );
  NAND2X1 U244 ( .A(N324), .B(n282), .Y(n285) );
  AOI22X1 U245 ( .A(N219), .B(n283), .C(X0[6]), .D(n606), .Y(n284) );
  NAND3X1 U246 ( .A(n287), .B(n288), .C(n289), .Y(n501) );
  AOI22X1 U247 ( .A(N331), .B(n280), .C(N210), .D(n281), .Y(n289) );
  NAND2X1 U248 ( .A(N323), .B(n282), .Y(n288) );
  AOI22X1 U249 ( .A(N218), .B(n283), .C(X0[5]), .D(n606), .Y(n287) );
  NAND3X1 U250 ( .A(n290), .B(n291), .C(n292), .Y(n502) );
  AOI22X1 U251 ( .A(N330), .B(n280), .C(N209), .D(n281), .Y(n292) );
  NAND2X1 U252 ( .A(N322), .B(n282), .Y(n291) );
  AOI22X1 U253 ( .A(N217), .B(n283), .C(X0[4]), .D(n606), .Y(n290) );
  OAI21X1 U254 ( .A(n576), .B(n629), .C(n293), .Y(n503) );
  AOI22X1 U255 ( .A(N232), .B(n9), .C(N216), .D(n1), .Y(n293) );
  OAI21X1 U256 ( .A(n576), .B(n628), .C(n294), .Y(n504) );
  AOI22X1 U257 ( .A(N231), .B(n9), .C(N215), .D(n1), .Y(n294) );
  OAI21X1 U258 ( .A(n576), .B(n627), .C(n295), .Y(n505) );
  AOI22X1 U259 ( .A(N230), .B(n9), .C(N214), .D(n1), .Y(n295) );
  OAI21X1 U260 ( .A(n576), .B(n642), .C(n296), .Y(n506) );
  AOI22X1 U261 ( .A(N229), .B(n9), .C(N213), .D(n1), .Y(n296) );
  NAND3X1 U263 ( .A(n298), .B(n235), .C(n577), .Y(n297) );
  NAND3X1 U264 ( .A(n299), .B(n300), .C(n301), .Y(n507) );
  AOI22X1 U265 ( .A(N329), .B(n280), .C(N232), .D(n281), .Y(n301) );
  NAND2X1 U266 ( .A(N321), .B(n282), .Y(n300) );
  AOI22X1 U267 ( .A(N216), .B(n283), .C(X0[3]), .D(n606), .Y(n299) );
  NAND3X1 U268 ( .A(n302), .B(n303), .C(n304), .Y(n508) );
  AOI22X1 U269 ( .A(N328), .B(n280), .C(N231), .D(n281), .Y(n304) );
  NAND2X1 U270 ( .A(N320), .B(n282), .Y(n303) );
  AOI22X1 U271 ( .A(N215), .B(n283), .C(X0[2]), .D(n606), .Y(n302) );
  NAND3X1 U272 ( .A(n305), .B(n306), .C(n307), .Y(n509) );
  AOI22X1 U273 ( .A(N327), .B(n280), .C(N230), .D(n281), .Y(n307) );
  NAND2X1 U274 ( .A(N319), .B(n282), .Y(n306) );
  AOI22X1 U275 ( .A(N214), .B(n283), .C(X0[1]), .D(n606), .Y(n305) );
  NAND3X1 U276 ( .A(n308), .B(n309), .C(n310), .Y(n510) );
  AOI22X1 U277 ( .A(N326), .B(n280), .C(N229), .D(n281), .Y(n310) );
  NOR2X1 U278 ( .A(n624), .B(n311), .Y(n280) );
  NAND2X1 U279 ( .A(N318), .B(n282), .Y(n309) );
  NOR2X1 U280 ( .A(n311), .B(iX), .Y(n282) );
  AOI22X1 U281 ( .A(N213), .B(n283), .C(X0[0]), .D(n606), .Y(n308) );
  NOR2X1 U282 ( .A(n281), .B(n243), .Y(n283) );
  NAND3X1 U283 ( .A(n313), .B(n314), .C(n315), .Y(n511) );
  AOI22X1 U284 ( .A(N296), .B(n316), .C(N220), .D(n317), .Y(n315) );
  NAND2X1 U285 ( .A(N288), .B(n318), .Y(n314) );
  AOI22X1 U286 ( .A(n319), .B(N212), .C(Y0[7]), .D(n606), .Y(n313) );
  NAND3X1 U287 ( .A(n320), .B(n321), .C(n322), .Y(n512) );
  AOI22X1 U288 ( .A(N295), .B(n316), .C(N219), .D(n317), .Y(n322) );
  NAND2X1 U289 ( .A(N287), .B(n318), .Y(n321) );
  AOI22X1 U290 ( .A(n319), .B(N211), .C(Y0[6]), .D(n606), .Y(n320) );
  NAND3X1 U291 ( .A(n323), .B(n324), .C(n325), .Y(n513) );
  AOI22X1 U292 ( .A(N294), .B(n316), .C(N218), .D(n317), .Y(n325) );
  NAND2X1 U293 ( .A(N286), .B(n318), .Y(n324) );
  AOI22X1 U294 ( .A(n319), .B(N210), .C(Y0[5]), .D(n606), .Y(n323) );
  NAND3X1 U295 ( .A(n326), .B(n327), .C(n328), .Y(n514) );
  AOI22X1 U296 ( .A(N293), .B(n316), .C(N217), .D(n317), .Y(n328) );
  NAND2X1 U297 ( .A(N285), .B(n318), .Y(n327) );
  AOI22X1 U298 ( .A(n319), .B(N209), .C(Y0[4]), .D(n606), .Y(n326) );
  NAND3X1 U299 ( .A(n329), .B(n330), .C(n331), .Y(n515) );
  AOI22X1 U300 ( .A(N292), .B(n316), .C(N216), .D(n317), .Y(n331) );
  NAND2X1 U301 ( .A(N284), .B(n318), .Y(n330) );
  AOI22X1 U302 ( .A(n319), .B(N232), .C(Y0[3]), .D(n606), .Y(n329) );
  NAND3X1 U303 ( .A(n332), .B(n333), .C(n334), .Y(n516) );
  AOI22X1 U304 ( .A(N291), .B(n316), .C(N215), .D(n317), .Y(n334) );
  NAND2X1 U305 ( .A(N283), .B(n318), .Y(n333) );
  AOI22X1 U306 ( .A(n319), .B(N231), .C(Y0[2]), .D(n606), .Y(n332) );
  NAND3X1 U307 ( .A(n335), .B(n336), .C(n337), .Y(n517) );
  AOI22X1 U308 ( .A(N290), .B(n316), .C(N214), .D(n317), .Y(n337) );
  NAND2X1 U309 ( .A(N282), .B(n318), .Y(n336) );
  AOI22X1 U310 ( .A(n319), .B(N230), .C(Y0[1]), .D(n606), .Y(n335) );
  NAND3X1 U311 ( .A(n338), .B(n339), .C(n340), .Y(n518) );
  AOI22X1 U312 ( .A(N289), .B(n316), .C(N213), .D(n317), .Y(n340) );
  NOR2X1 U313 ( .A(n625), .B(n341), .Y(n316) );
  NAND2X1 U314 ( .A(N281), .B(n318), .Y(n339) );
  NOR2X1 U315 ( .A(n341), .B(iY), .Y(n318) );
  AOI22X1 U316 ( .A(n319), .B(N229), .C(Y0[0]), .D(n606), .Y(n338) );
  NOR2X1 U317 ( .A(n317), .B(n243), .Y(n319) );
  NAND3X1 U318 ( .A(n342), .B(n298), .C(n343), .Y(n312) );
  NOR2X1 U319 ( .A(n607), .B(n605), .Y(n343) );
  OAI21X1 U320 ( .A(n594), .B(n624), .C(n344), .Y(n519) );
  OAI21X1 U321 ( .A(n345), .B(n346), .C(n594), .Y(n344) );
  OAI21X1 U323 ( .A(n594), .B(n625), .C(n347), .Y(n520) );
  OAI21X1 U324 ( .A(n348), .B(n349), .C(n594), .Y(n347) );
  NAND3X1 U326 ( .A(n254), .B(n242), .C(n342), .Y(n350) );
  AOI22X1 U327 ( .A(N264), .B(n601), .C(i[7]), .D(n352), .Y(n351) );
  AOI22X1 U328 ( .A(N263), .B(n601), .C(i[6]), .D(n352), .Y(n353) );
  AOI22X1 U329 ( .A(N262), .B(n601), .C(i[5]), .D(n352), .Y(n354) );
  AOI22X1 U330 ( .A(N261), .B(n601), .C(i[4]), .D(n352), .Y(n355) );
  AOI22X1 U331 ( .A(N260), .B(n601), .C(i[3]), .D(n352), .Y(n356) );
  AOI22X1 U332 ( .A(N259), .B(n601), .C(i[2]), .D(n352), .Y(n357) );
  AOI22X1 U333 ( .A(N258), .B(n601), .C(i[1]), .D(n352), .Y(n358) );
  NAND2X1 U334 ( .A(n359), .B(n360), .Y(n521) );
  AOI22X1 U336 ( .A(dy[8]), .B(n8), .C(dx[8]), .D(n7), .Y(n359) );
  NAND3X1 U337 ( .A(n364), .B(n365), .C(n366), .Y(n522) );
  AOI21X1 U338 ( .A(n10), .B(n7), .C(n593), .Y(n366) );
  AOI22X1 U339 ( .A(n8), .B(dy[7]), .C(n607), .D(n11), .Y(n367) );
  NAND2X1 U340 ( .A(N104), .B(n345), .Y(n365) );
  NAND3X1 U342 ( .A(n369), .B(n370), .C(n371), .Y(n523) );
  AOI21X1 U343 ( .A(n11), .B(n7), .C(n592), .Y(n371) );
  AOI22X1 U344 ( .A(n8), .B(dy[6]), .C(n607), .D(n12), .Y(n372) );
  NAND2X1 U345 ( .A(N103), .B(n345), .Y(n370) );
  NAND3X1 U347 ( .A(n373), .B(n374), .C(n375), .Y(n524) );
  AOI21X1 U348 ( .A(n12), .B(n7), .C(n591), .Y(n375) );
  AOI22X1 U349 ( .A(n8), .B(dy[5]), .C(n607), .D(n15), .Y(n376) );
  NAND2X1 U350 ( .A(N102), .B(n345), .Y(n374) );
  NAND3X1 U352 ( .A(n377), .B(n378), .C(n379), .Y(n525) );
  AOI21X1 U353 ( .A(n15), .B(n7), .C(n590), .Y(n379) );
  AOI22X1 U354 ( .A(n8), .B(dy[4]), .C(n607), .D(n18), .Y(n380) );
  NAND2X1 U355 ( .A(N101), .B(n345), .Y(n378) );
  NAND3X1 U357 ( .A(n381), .B(n382), .C(n383), .Y(n526) );
  AOI21X1 U358 ( .A(n18), .B(n7), .C(n589), .Y(n383) );
  AOI22X1 U359 ( .A(n8), .B(dy[3]), .C(n607), .D(n19), .Y(n384) );
  NAND2X1 U360 ( .A(N100), .B(n345), .Y(n382) );
  NAND3X1 U362 ( .A(n385), .B(n386), .C(n387), .Y(n527) );
  AOI21X1 U363 ( .A(n19), .B(n7), .C(n588), .Y(n387) );
  AOI22X1 U364 ( .A(n8), .B(dy[2]), .C(n607), .D(N190), .Y(n388) );
  NAND2X1 U365 ( .A(N99), .B(n345), .Y(n386) );
  NAND3X1 U367 ( .A(n389), .B(n390), .C(n391), .Y(n528) );
  AOI21X1 U368 ( .A(N190), .B(n7), .C(n587), .Y(n391) );
  AOI22X1 U369 ( .A(n8), .B(dy[1]), .C(n607), .D(dx[0]), .Y(n392) );
  NAND2X1 U370 ( .A(N98), .B(n345), .Y(n390) );
  NAND3X1 U372 ( .A(n393), .B(n394), .C(n395), .Y(n529) );
  AOI22X1 U373 ( .A(dy[0]), .B(n8), .C(dx[0]), .D(n7), .Y(n395) );
  NAND2X1 U375 ( .A(N97), .B(n345), .Y(n394) );
  NOR2X1 U376 ( .A(n566), .B(n262), .Y(n345) );
  NOR2X1 U378 ( .A(n262), .B(N95), .Y(n368) );
  NAND2X1 U380 ( .A(n396), .B(n397), .Y(n530) );
  AOI22X1 U382 ( .A(dx[8]), .B(n8), .C(dy[8]), .D(n363), .Y(n396) );
  NAND3X1 U383 ( .A(n400), .B(n401), .C(n402), .Y(n531) );
  AOI21X1 U384 ( .A(dy[7]), .B(n363), .C(n586), .Y(n402) );
  AOI22X1 U385 ( .A(n10), .B(n8), .C(n607), .D(dy[6]), .Y(n403) );
  NAND2X1 U386 ( .A(N130), .B(n348), .Y(n401) );
  NAND3X1 U388 ( .A(n405), .B(n406), .C(n407), .Y(n532) );
  AOI21X1 U389 ( .A(dy[6]), .B(n363), .C(n585), .Y(n407) );
  AOI22X1 U390 ( .A(n8), .B(n11), .C(n607), .D(dy[5]), .Y(n408) );
  NAND2X1 U391 ( .A(N129), .B(n348), .Y(n406) );
  NAND3X1 U393 ( .A(n409), .B(n410), .C(n411), .Y(n533) );
  AOI21X1 U394 ( .A(dy[5]), .B(n363), .C(n584), .Y(n411) );
  AOI22X1 U395 ( .A(n8), .B(n12), .C(n607), .D(dy[4]), .Y(n412) );
  NAND2X1 U396 ( .A(N128), .B(n348), .Y(n410) );
  NAND3X1 U398 ( .A(n413), .B(n414), .C(n415), .Y(n534) );
  AOI21X1 U399 ( .A(dy[4]), .B(n363), .C(n583), .Y(n415) );
  AOI22X1 U400 ( .A(n8), .B(n15), .C(n607), .D(dy[3]), .Y(n416) );
  NAND2X1 U401 ( .A(N127), .B(n348), .Y(n414) );
  NAND3X1 U403 ( .A(n417), .B(n418), .C(n419), .Y(n535) );
  AOI21X1 U404 ( .A(dy[3]), .B(n363), .C(n582), .Y(n419) );
  AOI22X1 U405 ( .A(n8), .B(n18), .C(n607), .D(dy[2]), .Y(n420) );
  NAND2X1 U406 ( .A(N126), .B(n348), .Y(n418) );
  NAND3X1 U408 ( .A(n421), .B(n422), .C(n423), .Y(n536) );
  AOI21X1 U409 ( .A(dy[2]), .B(n363), .C(n581), .Y(n423) );
  AOI22X1 U410 ( .A(n8), .B(n19), .C(n607), .D(dy[1]), .Y(n424) );
  NAND2X1 U411 ( .A(N125), .B(n348), .Y(n422) );
  NAND3X1 U413 ( .A(n425), .B(n426), .C(n427), .Y(n537) );
  AOI21X1 U414 ( .A(dy[1]), .B(n363), .C(n580), .Y(n427) );
  AOI22X1 U415 ( .A(n8), .B(N190), .C(n607), .D(dy[0]), .Y(n428) );
  NAND2X1 U416 ( .A(N124), .B(n348), .Y(n426) );
  NAND3X1 U418 ( .A(n429), .B(n430), .C(n431), .Y(n538) );
  AOI22X1 U419 ( .A(dx[0]), .B(n8), .C(dy[0]), .D(n363), .Y(n431) );
  NAND3X1 U422 ( .A(n254), .B(n298), .C(n342), .Y(n432) );
  NOR3X1 U423 ( .A(n603), .B(n609), .C(n433), .Y(n342) );
  OAI21X1 U424 ( .A(n243), .B(steep), .C(n595), .Y(n433) );
  NAND2X1 U425 ( .A(N123), .B(n348), .Y(n430) );
  NOR2X1 U426 ( .A(n565), .B(n262), .Y(n348) );
  NOR2X1 U428 ( .A(n262), .B(N121), .Y(n404) );
  OAI21X1 U430 ( .A(n242), .B(n613), .C(n434), .Y(n539) );
  OAI21X1 U431 ( .A(n602), .B(n435), .C(steep), .Y(n434) );
  NAND2X1 U432 ( .A(n437), .B(n438), .Y(n540) );
  AOI22X1 U433 ( .A(N199), .B(n603), .C(N306), .D(n611), .Y(n438) );
  AOI22X1 U434 ( .A(N269), .B(n612), .C(err[0]), .D(n578), .Y(n437) );
  NAND2X1 U435 ( .A(n439), .B(n440), .Y(n541) );
  AOI22X1 U436 ( .A(N200), .B(n603), .C(N307), .D(n611), .Y(n440) );
  AOI22X1 U437 ( .A(N270), .B(n612), .C(err[1]), .D(n578), .Y(n439) );
  NAND2X1 U438 ( .A(n441), .B(n442), .Y(n542) );
  AOI22X1 U439 ( .A(N201), .B(n603), .C(N308), .D(n611), .Y(n442) );
  AOI22X1 U440 ( .A(N271), .B(n612), .C(err[2]), .D(n578), .Y(n441) );
  NAND2X1 U441 ( .A(n443), .B(n444), .Y(n543) );
  AOI22X1 U442 ( .A(N202), .B(n603), .C(N309), .D(n611), .Y(n444) );
  AOI22X1 U443 ( .A(N272), .B(n612), .C(err[3]), .D(n578), .Y(n443) );
  NAND2X1 U444 ( .A(n445), .B(n446), .Y(n544) );
  AOI22X1 U445 ( .A(N203), .B(n603), .C(N310), .D(n611), .Y(n446) );
  AOI22X1 U446 ( .A(N273), .B(n612), .C(err[4]), .D(n578), .Y(n445) );
  NAND2X1 U447 ( .A(n447), .B(n448), .Y(n545) );
  AOI22X1 U448 ( .A(N204), .B(n603), .C(N311), .D(n611), .Y(n448) );
  AOI22X1 U449 ( .A(N274), .B(n612), .C(err[5]), .D(n578), .Y(n447) );
  NAND2X1 U450 ( .A(n449), .B(n450), .Y(n546) );
  AOI22X1 U451 ( .A(N205), .B(n603), .C(N312), .D(n611), .Y(n450) );
  AOI22X1 U452 ( .A(N275), .B(n612), .C(err[6]), .D(n578), .Y(n449) );
  NAND2X1 U453 ( .A(n451), .B(n452), .Y(n547) );
  AOI22X1 U454 ( .A(N206), .B(n603), .C(N313), .D(n611), .Y(n452) );
  AOI22X1 U455 ( .A(N276), .B(n612), .C(err[7]), .D(n578), .Y(n451) );
  OAI21X1 U456 ( .A(n453), .B(n626), .C(n454), .Y(n548) );
  AOI22X1 U457 ( .A(N315), .B(n611), .C(N278), .D(n612), .Y(n454) );
  OAI21X1 U458 ( .A(n453), .B(n615), .C(n455), .Y(n549) );
  AOI22X1 U459 ( .A(N316), .B(n611), .C(N279), .D(n612), .Y(n455) );
  OAI22X1 U460 ( .A(n600), .B(n618), .C(n456), .D(n457), .Y(n550) );
  XNOR2X1 U461 ( .A(count[3]), .B(n458), .Y(n457) );
  NOR2X1 U462 ( .A(n623), .B(n620), .Y(n458) );
  OAI21X1 U463 ( .A(n459), .B(n623), .C(n460), .Y(n551) );
  NAND3X1 U464 ( .A(n575), .B(n623), .C(n461), .Y(n460) );
  AOI21X1 U465 ( .A(n620), .B(n575), .C(n462), .Y(n459) );
  NOR2X1 U466 ( .A(n622), .B(n621), .Y(n461) );
  OAI21X1 U467 ( .A(n463), .B(n622), .C(n464), .Y(n552) );
  NAND3X1 U468 ( .A(n575), .B(n622), .C(count[0]), .Y(n464) );
  AOI21X1 U469 ( .A(n575), .B(n621), .C(n462), .Y(n463) );
  OAI22X1 U470 ( .A(n600), .B(n621), .C(count[0]), .D(n456), .Y(n553) );
  NAND3X1 U471 ( .A(n436), .B(n465), .C(n466), .Y(n462) );
  NOR2X1 U472 ( .A(n608), .B(n467), .Y(n466) );
  NAND2X1 U473 ( .A(n256), .B(n242), .Y(n467) );
  OAI21X1 U474 ( .A(n453), .B(n614), .C(n468), .Y(n554) );
  AOI22X1 U475 ( .A(N317), .B(n611), .C(N280), .D(n612), .Y(n468) );
  NAND3X1 U476 ( .A(n469), .B(n470), .C(n471), .Y(n555) );
  AOI21X1 U477 ( .A(err[8]), .B(n578), .C(n608), .Y(n471) );
  NAND2X1 U478 ( .A(n472), .B(n473), .Y(n298) );
  NOR2X1 U479 ( .A(n474), .B(n475), .Y(n453) );
  NAND3X1 U480 ( .A(n255), .B(n262), .C(n595), .Y(n475) );
  NAND3X1 U481 ( .A(n248), .B(n235), .C(n596), .Y(n435) );
  NAND3X1 U482 ( .A(n243), .B(n234), .C(n242), .Y(n474) );
  NAND2X1 U483 ( .A(N277), .B(n612), .Y(n470) );
  AOI22X1 U484 ( .A(N207), .B(n603), .C(N314), .D(n611), .Y(n469) );
  AOI22X1 U485 ( .A(N257), .B(n601), .C(i[0]), .D(n352), .Y(n476) );
  NAND2X1 U486 ( .A(n577), .B(n248), .Y(n352) );
  NAND2X1 U487 ( .A(n477), .B(n478), .Y(n248) );
  NAND3X1 U488 ( .A(n436), .B(n242), .C(n596), .Y(n479) );
  NAND3X1 U489 ( .A(n256), .B(n456), .C(n465), .Y(n480) );
  NAND2X1 U490 ( .A(state[1]), .B(n481), .Y(n465) );
  NOR2X1 U491 ( .A(rast_done), .B(n599), .Y(n456) );
  NAND2X1 U492 ( .A(n481), .B(n482), .Y(n244) );
  NAND2X1 U493 ( .A(n483), .B(n484), .Y(n256) );
  NAND2X1 U494 ( .A(n472), .B(n484), .Y(n242) );
  NOR2X1 U495 ( .A(n485), .B(n486), .Y(n436) );
  NAND3X1 U496 ( .A(n255), .B(n262), .C(n254), .Y(n486) );
  NOR2X1 U497 ( .A(n611), .B(n612), .Y(n254) );
  NAND2X1 U498 ( .A(n483), .B(n482), .Y(n341) );
  NAND2X1 U499 ( .A(n477), .B(n483), .Y(n311) );
  NAND2X1 U500 ( .A(n472), .B(n482), .Y(n262) );
  NAND2X1 U501 ( .A(n472), .B(n477), .Y(n255) );
  NOR2X1 U502 ( .A(state[2]), .B(state[3]), .Y(n472) );
  NAND3X1 U503 ( .A(n243), .B(n234), .C(n241), .Y(n485) );
  NAND2X1 U504 ( .A(n478), .B(n482), .Y(n241) );
  NOR2X1 U505 ( .A(n616), .B(state[1]), .Y(n482) );
  NAND2X1 U506 ( .A(n473), .B(n483), .Y(n234) );
  NOR2X1 U507 ( .A(n619), .B(state[2]), .Y(n483) );
  NAND2X1 U508 ( .A(n473), .B(n478), .Y(n243) );
  NAND2X1 U509 ( .A(n478), .B(n484), .Y(n235) );
  NOR2X1 U510 ( .A(n604), .B(state[3]), .Y(n478) );
  NAND2X1 U511 ( .A(n473), .B(n481), .Y(n247) );
  NOR2X1 U512 ( .A(n619), .B(n604), .Y(n481) );
  NOR2X1 U513 ( .A(state[0]), .B(state[1]), .Y(n473) );
  Rasterizer_DW01_inc_0 add_262 ( .A({N212, N211, N210, N209, N232, N231, N230, 
        N229}), .SUM({N325, N324, N323, N322, N321, N320, N319, N318}) );
  Rasterizer_DW01_add_0 add_259 ( .A(err), .B({1'b0, 1'b0, 1'b0, dy}), .CI(
        1'b0), .SUM({N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307, N306}) );
  Rasterizer_DW01_inc_1 add_249 ( .A({N220, N219, N218, N217, N216, N215, N214, 
        N213}), .SUM({N288, N287, N286, N285, N284, N283, N282, N281}) );
  Rasterizer_DW01_sub_2 sub_246 ( .A(err), .B({1'b0, 1'b0, 1'b0, dx[8], n10, 
        n11, n12, n15, n18, n19, N190, dx[0]}), .CI(1'b0), .DIFF({N280, N279, 
        N278, N277, N276, N275, N274, N273, N272, N271, N270, N269}) );
  Rasterizer_DW01_inc_2 add_222 ( .A(i), .SUM({N264, N263, N262, N261, N260, 
        N259, N258, N257}) );
  Rasterizer_DW01_sub_3 sub_126 ( .A(Y1), .B(Y0), .CI(1'b0), .DIFF({N138, N137, 
        N136, N135, N134, N133, N132, N131}) );
  Rasterizer_DW01_sub_4 sub_123 ( .A(Y0), .B(Y1), .CI(1'b0), .DIFF({N130, N129, 
        N128, N127, N126, N125, N124, N123}) );
  Rasterizer_DW01_sub_5 sub_116 ( .A(X1), .B(X0), .CI(1'b0), .DIFF({N112, N111, 
        N110, N109, N108, N107, N106, N105}) );
  Rasterizer_DW01_sub_6 sub_111 ( .A(X0), .B(X1), .CI(1'b0), .DIFF({N104, N103, 
        N102, N101, N100, N99, N98, N97}) );
  Rasterizer_DW01_add_3 add_0_root_sub_0_root_sub_184 ( .A(dy), .B({N198, N197, 
        N196, N195, N194, N193, N192, N191, N190}), .CI(1'b0), .SUM({N207, 
        N206, N205, N204, N203, N202, N201, N200, N199}) );
  AND2X2 U13 ( .A(steep), .B(n576), .Y(n1) );
  INVX2 U14 ( .A(n297), .Y(n576) );
  INVX2 U17 ( .A(n2), .Y(n8) );
  INVX2 U18 ( .A(n453), .Y(n578) );
  OR2X2 U19 ( .A(n432), .B(n243), .Y(n2) );
  INVX2 U20 ( .A(n311), .Y(n611) );
  INVX2 U21 ( .A(n341), .Y(n612) );
  INVX2 U22 ( .A(n6), .Y(n7) );
  INVX2 U23 ( .A(n363), .Y(n6) );
  INVX2 U24 ( .A(n242), .Y(n607) );
  INVX2 U27 ( .A(n241), .Y(n603) );
  INVX2 U30 ( .A(n262), .Y(n606) );
  INVX2 U103 ( .A(n235), .Y(n601) );
  INVX2 U108 ( .A(n5), .Y(n9) );
  BUFX2 U109 ( .A(dx[2]), .Y(n19) );
  BUFX2 U110 ( .A(dx[3]), .Y(n18) );
  INVX2 U111 ( .A(N190), .Y(n20) );
  OR2X2 U112 ( .A(n297), .B(steep), .Y(n5) );
  BUFX2 U113 ( .A(dx[5]), .Y(n12) );
  BUFX2 U114 ( .A(dx[4]), .Y(n15) );
  BUFX2 U115 ( .A(dx[6]), .Y(n11) );
  BUFX2 U116 ( .A(dx[7]), .Y(n10) );
  BUFX2 U117 ( .A(RST_N), .Y(n26) );
  BUFX2 U118 ( .A(RST_N), .Y(n25) );
  BUFX2 U119 ( .A(RST_N), .Y(n23) );
  BUFX2 U120 ( .A(RST_N), .Y(n22) );
  BUFX2 U121 ( .A(RST_N), .Y(n21) );
  BUFX2 U122 ( .A(RST_N), .Y(n24) );
  BUFX2 U123 ( .A(RST_N), .Y(n27) );
  INVX1 U124 ( .A(Y1[7]), .Y(n195) );
  AND2X1 U125 ( .A(n28), .B(\sub_1_root_sub_0_root_sub_184/carry[7] ), .Y(N198) );
  XOR2X1 U126 ( .A(\sub_1_root_sub_0_root_sub_184/carry[7] ), .B(n28), .Y(N197) );
  AND2X1 U127 ( .A(n29), .B(\sub_1_root_sub_0_root_sub_184/carry[6] ), .Y(
        \sub_1_root_sub_0_root_sub_184/carry[7] ) );
  XOR2X1 U128 ( .A(\sub_1_root_sub_0_root_sub_184/carry[6] ), .B(n29), .Y(N196) );
  AND2X1 U129 ( .A(n30), .B(\sub_1_root_sub_0_root_sub_184/carry[5] ), .Y(
        \sub_1_root_sub_0_root_sub_184/carry[6] ) );
  XOR2X1 U130 ( .A(\sub_1_root_sub_0_root_sub_184/carry[5] ), .B(n30), .Y(N195) );
  AND2X1 U131 ( .A(n31), .B(\sub_1_root_sub_0_root_sub_184/carry[4] ), .Y(
        \sub_1_root_sub_0_root_sub_184/carry[5] ) );
  XOR2X1 U132 ( .A(\sub_1_root_sub_0_root_sub_184/carry[4] ), .B(n31), .Y(N194) );
  AND2X1 U133 ( .A(n32), .B(\sub_1_root_sub_0_root_sub_184/carry[3] ), .Y(
        \sub_1_root_sub_0_root_sub_184/carry[4] ) );
  XOR2X1 U134 ( .A(\sub_1_root_sub_0_root_sub_184/carry[3] ), .B(n32), .Y(N193) );
  AND2X1 U135 ( .A(n33), .B(\sub_1_root_sub_0_root_sub_184/carry[2] ), .Y(
        \sub_1_root_sub_0_root_sub_184/carry[3] ) );
  XOR2X1 U136 ( .A(\sub_1_root_sub_0_root_sub_184/carry[2] ), .B(n33), .Y(N192) );
  AND2X1 U137 ( .A(n34), .B(n20), .Y(\sub_1_root_sub_0_root_sub_184/carry[2] )
         );
  XOR2X1 U138 ( .A(n20), .B(n34), .Y(N191) );
  INVX2 U139 ( .A(dx[8]), .Y(n28) );
  INVX2 U140 ( .A(n10), .Y(n29) );
  INVX2 U141 ( .A(n11), .Y(n30) );
  INVX2 U142 ( .A(n12), .Y(n31) );
  INVX2 U143 ( .A(n15), .Y(n32) );
  INVX2 U144 ( .A(n18), .Y(n33) );
  INVX2 U145 ( .A(n19), .Y(n34) );
  NAND2X1 U146 ( .A(n44), .B(N289), .Y(n35) );
  OAI21X1 U147 ( .A(N289), .B(n44), .C(n35), .Y(N290) );
  NOR2X1 U148 ( .A(n35), .B(N215), .Y(n37) );
  AOI21X1 U149 ( .A(n35), .B(N215), .C(n37), .Y(n36) );
  NAND2X1 U150 ( .A(n37), .B(n43), .Y(n38) );
  OAI21X1 U151 ( .A(n37), .B(n43), .C(n38), .Y(N292) );
  NOR2X1 U152 ( .A(n38), .B(N217), .Y(n40) );
  AOI21X1 U153 ( .A(n38), .B(N217), .C(n40), .Y(n39) );
  NAND2X1 U154 ( .A(n40), .B(n45), .Y(n41) );
  OAI21X1 U155 ( .A(n40), .B(n45), .C(n41), .Y(N294) );
  XNOR2X1 U156 ( .A(N219), .B(n41), .Y(N295) );
  NOR2X1 U157 ( .A(N219), .B(n41), .Y(n42) );
  XOR2X1 U158 ( .A(N220), .B(n42), .Y(N296) );
  INVX2 U159 ( .A(N216), .Y(n43) );
  INVX2 U160 ( .A(N214), .Y(n44) );
  INVX2 U161 ( .A(N218), .Y(n45) );
  INVX2 U162 ( .A(N213), .Y(N289) );
  INVX2 U163 ( .A(n39), .Y(N293) );
  INVX2 U164 ( .A(n36), .Y(N291) );
  NAND2X1 U165 ( .A(n55), .B(N326), .Y(n46) );
  OAI21X1 U166 ( .A(N326), .B(n55), .C(n46), .Y(N327) );
  NOR2X1 U167 ( .A(n46), .B(N231), .Y(n48) );
  AOI21X1 U168 ( .A(n46), .B(N231), .C(n48), .Y(n47) );
  NAND2X1 U169 ( .A(n48), .B(n54), .Y(n49) );
  OAI21X1 U170 ( .A(n48), .B(n54), .C(n49), .Y(N329) );
  NOR2X1 U171 ( .A(n49), .B(N209), .Y(n51) );
  AOI21X1 U172 ( .A(n49), .B(N209), .C(n51), .Y(n50) );
  NAND2X1 U173 ( .A(n51), .B(n56), .Y(n52) );
  OAI21X1 U174 ( .A(n51), .B(n56), .C(n52), .Y(N331) );
  XNOR2X1 U175 ( .A(N211), .B(n52), .Y(N332) );
  NOR2X1 U176 ( .A(N211), .B(n52), .Y(n53) );
  XOR2X1 U177 ( .A(N212), .B(n53), .Y(N333) );
  INVX2 U178 ( .A(N232), .Y(n54) );
  INVX2 U179 ( .A(N230), .Y(n55) );
  INVX2 U180 ( .A(N210), .Y(n56) );
  INVX2 U181 ( .A(N229), .Y(N326) );
  INVX2 U182 ( .A(n50), .Y(N330) );
  INVX2 U183 ( .A(n47), .Y(N328) );
  NAND2X1 U184 ( .A(X0[0]), .B(n152), .Y(n58) );
  OAI21X1 U185 ( .A(n58), .B(X1[1]), .C(n153), .Y(n57) );
  AOI21X1 U186 ( .A(X1[1]), .B(n58), .C(n154), .Y(n59) );
  OAI21X1 U187 ( .A(X0[2]), .B(n156), .C(n59), .Y(n60) );
  OAI21X1 U262 ( .A(X1[2]), .B(n155), .C(n60), .Y(n61) );
  AOI21X1 U322 ( .A(X0[3]), .B(n158), .C(n61), .Y(n62) );
  AOI21X1 U325 ( .A(X1[3]), .B(n157), .C(n62), .Y(n63) );
  OAI21X1 U335 ( .A(X0[4]), .B(n160), .C(n63), .Y(n64) );
  OAI21X1 U341 ( .A(X1[4]), .B(n159), .C(n64), .Y(n65) );
  AOI21X1 U346 ( .A(X0[5]), .B(n162), .C(n65), .Y(n66) );
  AOI21X1 U351 ( .A(X1[5]), .B(n161), .C(n66), .Y(n67) );
  OAI21X1 U356 ( .A(X0[6]), .B(n164), .C(n67), .Y(n149) );
  OAI21X1 U361 ( .A(X1[6]), .B(n163), .C(n149), .Y(n150) );
  OAI21X1 U366 ( .A(X0[7]), .B(n166), .C(n150), .Y(n151) );
  OAI21X1 U371 ( .A(X1[7]), .B(n165), .C(n151), .Y(N95) );
  INVX2 U374 ( .A(X1[0]), .Y(n152) );
  INVX2 U377 ( .A(X0[1]), .Y(n153) );
  INVX2 U379 ( .A(n57), .Y(n154) );
  INVX2 U381 ( .A(X0[2]), .Y(n155) );
  INVX2 U387 ( .A(X1[2]), .Y(n156) );
  INVX2 U392 ( .A(X0[3]), .Y(n157) );
  INVX2 U397 ( .A(X1[3]), .Y(n158) );
  INVX2 U402 ( .A(X0[4]), .Y(n159) );
  INVX2 U407 ( .A(X1[4]), .Y(n160) );
  INVX2 U412 ( .A(X0[5]), .Y(n161) );
  INVX2 U417 ( .A(X1[5]), .Y(n162) );
  INVX2 U420 ( .A(X0[6]), .Y(n163) );
  INVX2 U421 ( .A(X1[6]), .Y(n164) );
  INVX2 U427 ( .A(X0[7]), .Y(n165) );
  INVX2 U429 ( .A(X1[7]), .Y(n166) );
  NAND2X1 U514 ( .A(Y0[0]), .B(n181), .Y(n168) );
  OAI21X1 U515 ( .A(n168), .B(Y1[1]), .C(n182), .Y(n167) );
  AOI21X1 U516 ( .A(Y1[1]), .B(n168), .C(n183), .Y(n169) );
  OAI21X1 U517 ( .A(Y0[2]), .B(n185), .C(n169), .Y(n170) );
  OAI21X1 U518 ( .A(Y1[2]), .B(n184), .C(n170), .Y(n171) );
  AOI21X1 U519 ( .A(Y0[3]), .B(n187), .C(n171), .Y(n172) );
  AOI21X1 U520 ( .A(Y1[3]), .B(n186), .C(n172), .Y(n173) );
  OAI21X1 U521 ( .A(Y0[4]), .B(n189), .C(n173), .Y(n174) );
  OAI21X1 U522 ( .A(Y1[4]), .B(n188), .C(n174), .Y(n175) );
  AOI21X1 U523 ( .A(Y0[5]), .B(n191), .C(n175), .Y(n176) );
  AOI21X1 U524 ( .A(Y1[5]), .B(n190), .C(n176), .Y(n177) );
  OAI21X1 U525 ( .A(Y0[6]), .B(n193), .C(n177), .Y(n178) );
  OAI21X1 U526 ( .A(Y1[6]), .B(n192), .C(n178), .Y(n179) );
  OAI21X1 U527 ( .A(Y0[7]), .B(n195), .C(n179), .Y(n180) );
  OAI21X1 U528 ( .A(Y1[7]), .B(n194), .C(n180), .Y(N121) );
  INVX2 U529 ( .A(Y1[0]), .Y(n181) );
  INVX2 U530 ( .A(Y0[1]), .Y(n182) );
  INVX2 U531 ( .A(n167), .Y(n183) );
  INVX2 U532 ( .A(Y0[2]), .Y(n184) );
  INVX2 U533 ( .A(Y1[2]), .Y(n185) );
  INVX2 U534 ( .A(Y0[3]), .Y(n186) );
  INVX2 U535 ( .A(Y1[3]), .Y(n187) );
  INVX2 U536 ( .A(Y0[4]), .Y(n188) );
  INVX2 U537 ( .A(Y1[4]), .Y(n189) );
  INVX2 U538 ( .A(Y0[5]), .Y(n190) );
  INVX2 U539 ( .A(Y1[5]), .Y(n191) );
  INVX2 U540 ( .A(Y0[6]), .Y(n192) );
  INVX2 U541 ( .A(Y1[6]), .Y(n193) );
  INVX2 U542 ( .A(Y0[7]), .Y(n194) );
  NAND2X1 U543 ( .A(dy[0]), .B(n220), .Y(n197) );
  OAI21X1 U544 ( .A(n197), .B(N190), .C(n217), .Y(n196) );
  AOI21X1 U545 ( .A(N190), .B(n197), .C(n221), .Y(n198) );
  OAI21X1 U546 ( .A(dy[2]), .B(n34), .C(n198), .Y(n199) );
  OAI21X1 U547 ( .A(n19), .B(n216), .C(n199), .Y(n200) );
  AOI21X1 U548 ( .A(dy[3]), .B(n33), .C(n200), .Y(n201) );
  AOI21X1 U549 ( .A(n18), .B(n215), .C(n201), .Y(n202) );
  OAI21X1 U550 ( .A(dy[4]), .B(n32), .C(n202), .Y(n203) );
  OAI21X1 U551 ( .A(n15), .B(n214), .C(n203), .Y(n204) );
  AOI21X1 U552 ( .A(dy[5]), .B(n31), .C(n204), .Y(n205) );
  AOI21X1 U553 ( .A(n12), .B(n213), .C(n205), .Y(n206) );
  OAI21X1 U554 ( .A(dy[6]), .B(n30), .C(n206), .Y(n207) );
  OAI21X1 U555 ( .A(n11), .B(n212), .C(n207), .Y(n208) );
  AOI21X1 U556 ( .A(dy[7]), .B(n29), .C(n208), .Y(n209) );
  AOI21X1 U557 ( .A(n10), .B(n218), .C(n209), .Y(n210) );
  OAI21X1 U558 ( .A(dy[8]), .B(n28), .C(n210), .Y(n211) );
  OAI21X1 U559 ( .A(dx[8]), .B(n219), .C(n211), .Y(N188) );
  INVX2 U560 ( .A(dy[6]), .Y(n212) );
  INVX2 U561 ( .A(dy[5]), .Y(n213) );
  INVX2 U562 ( .A(dy[4]), .Y(n214) );
  INVX2 U563 ( .A(dy[3]), .Y(n215) );
  INVX2 U564 ( .A(dy[2]), .Y(n216) );
  INVX2 U565 ( .A(dy[1]), .Y(n217) );
  INVX2 U566 ( .A(dy[7]), .Y(n218) );
  INVX2 U567 ( .A(dy[8]), .Y(n219) );
  INVX2 U568 ( .A(dx[0]), .Y(n220) );
  INVX2 U569 ( .A(n196), .Y(n221) );
  AOI21X1 U570 ( .A(i[1]), .B(n34), .C(i[0]), .Y(n222) );
  AOI22X1 U571 ( .A(n222), .B(N190), .C(n19), .D(n561), .Y(n223) );
  OAI21X1 U572 ( .A(i[2]), .B(n33), .C(n223), .Y(n224) );
  OAI21X1 U573 ( .A(n18), .B(n560), .C(n224), .Y(n225) );
  AOI21X1 U574 ( .A(i[3]), .B(n32), .C(n225), .Y(n226) );
  AOI21X1 U575 ( .A(n15), .B(n559), .C(n226), .Y(n227) );
  OAI21X1 U576 ( .A(i[4]), .B(n31), .C(n227), .Y(n228) );
  OAI21X1 U577 ( .A(n12), .B(n558), .C(n228), .Y(n264) );
  AOI21X1 U578 ( .A(i[5]), .B(n30), .C(n264), .Y(n265) );
  AOI21X1 U579 ( .A(n11), .B(n557), .C(n265), .Y(n361) );
  OAI21X1 U580 ( .A(i[6]), .B(n29), .C(n361), .Y(n362) );
  OAI21X1 U581 ( .A(n10), .B(n556), .C(n362), .Y(n398) );
  OAI21X1 U582 ( .A(i[7]), .B(n28), .C(n398), .Y(n399) );
  OAI21X1 U583 ( .A(dx[8]), .B(n562), .C(n399), .Y(N265) );
  INVX2 U584 ( .A(i[6]), .Y(n556) );
  INVX2 U585 ( .A(i[5]), .Y(n557) );
  INVX2 U586 ( .A(i[4]), .Y(n558) );
  INVX2 U587 ( .A(i[3]), .Y(n559) );
  INVX2 U588 ( .A(i[2]), .Y(n560) );
  INVX2 U589 ( .A(i[1]), .Y(n561) );
  INVX2 U590 ( .A(i[7]), .Y(n562) );
  NOR2X1 U591 ( .A(err[11]), .B(err[10]), .Y(n564) );
  NOR2X1 U592 ( .A(err[9]), .B(err[8]), .Y(n563) );
  NAND2X1 U593 ( .A(n564), .B(n563), .Y(N266) );
  INVX2 U594 ( .A(N121), .Y(n565) );
  INVX2 U595 ( .A(N95), .Y(n566) );
  INVX2 U596 ( .A(n476), .Y(n567) );
  INVX2 U597 ( .A(n351), .Y(n568) );
  INVX2 U598 ( .A(n353), .Y(n569) );
  INVX2 U599 ( .A(n354), .Y(n570) );
  INVX2 U600 ( .A(n355), .Y(n571) );
  INVX2 U601 ( .A(n356), .Y(n572) );
  INVX2 U602 ( .A(n357), .Y(n573) );
  INVX2 U603 ( .A(n358), .Y(n574) );
  INVX2 U604 ( .A(n456), .Y(n575) );
  INVX2 U605 ( .A(n479), .Y(n577) );
  INVX2 U606 ( .A(n432), .Y(n579) );
  INVX2 U607 ( .A(n428), .Y(n580) );
  INVX2 U608 ( .A(n424), .Y(n581) );
  INVX2 U609 ( .A(n420), .Y(n582) );
  INVX2 U610 ( .A(n416), .Y(n583) );
  INVX2 U611 ( .A(n412), .Y(n584) );
  INVX2 U612 ( .A(n408), .Y(n585) );
  INVX2 U613 ( .A(n403), .Y(n586) );
  INVX2 U614 ( .A(n392), .Y(n587) );
  INVX2 U615 ( .A(n388), .Y(n588) );
  INVX2 U616 ( .A(n384), .Y(n589) );
  INVX2 U617 ( .A(n380), .Y(n590) );
  INVX2 U618 ( .A(n376), .Y(n591) );
  INVX2 U619 ( .A(n372), .Y(n592) );
  INVX2 U620 ( .A(n367), .Y(n593) );
  INVX2 U621 ( .A(n350), .Y(n594) );
  INVX2 U622 ( .A(n435), .Y(n595) );
  INVX2 U623 ( .A(n480), .Y(n596) );
  INVX2 U624 ( .A(n247), .Y(rast_done) );
  INVX2 U625 ( .A(n245), .Y(n598) );
  INVX2 U626 ( .A(n244), .Y(n599) );
  INVX2 U627 ( .A(n462), .Y(n600) );
  INVX2 U628 ( .A(n436), .Y(n602) );
  INVX2 U629 ( .A(state[2]), .Y(n604) );
  INVX2 U630 ( .A(n255), .Y(n605) );
  INVX2 U631 ( .A(n298), .Y(n608) );
  INVX2 U632 ( .A(n234), .Y(n609) );
  INVX2 U633 ( .A(n254), .Y(n610) );
  INVX2 U634 ( .A(N188), .Y(n613) );
  INVX2 U635 ( .A(err[11]), .Y(n614) );
  INVX2 U636 ( .A(err[10]), .Y(n615) );
  INVX2 U637 ( .A(state[0]), .Y(n616) );
  INVX2 U638 ( .A(n236), .Y(n617) );
  INVX2 U639 ( .A(count[3]), .Y(n618) );
  INVX2 U640 ( .A(state[3]), .Y(n619) );
  INVX2 U641 ( .A(n461), .Y(n620) );
  INVX2 U642 ( .A(count[0]), .Y(n621) );
  INVX2 U643 ( .A(count[1]), .Y(n622) );
  INVX2 U644 ( .A(count[2]), .Y(n623) );
  INVX2 U645 ( .A(iX), .Y(n624) );
  INVX2 U646 ( .A(iY), .Y(n625) );
  INVX2 U647 ( .A(err[9]), .Y(n626) );
  INVX2 U648 ( .A(rast_index[1]), .Y(n627) );
  INVX2 U649 ( .A(rast_index[2]), .Y(n628) );
  INVX2 U650 ( .A(rast_index[3]), .Y(n629) );
  INVX2 U651 ( .A(rast_addr[0]), .Y(n630) );
  INVX2 U652 ( .A(rast_addr[1]), .Y(n631) );
  INVX2 U653 ( .A(rast_addr[2]), .Y(n632) );
  INVX2 U654 ( .A(rast_addr[3]), .Y(n633) );
  INVX2 U655 ( .A(rast_addr[4]), .Y(n634) );
  INVX2 U656 ( .A(rast_addr[5]), .Y(n635) );
  INVX2 U657 ( .A(rast_addr[6]), .Y(n636) );
  INVX2 U658 ( .A(rast_addr[7]), .Y(n637) );
  INVX2 U659 ( .A(rast_addr[8]), .Y(n638) );
  INVX2 U660 ( .A(rast_addr[9]), .Y(n639) );
  INVX2 U661 ( .A(rast_addr[10]), .Y(n640) );
  INVX2 U662 ( .A(rast_addr[11]), .Y(n641) );
  INVX2 U663 ( .A(rast_index[0]), .Y(n642) );
  OAI21X1 U664 ( .A(n243), .B(n624), .C(n255), .Y(n349) );
  OAI21X1 U665 ( .A(n243), .B(n625), .C(n255), .Y(n346) );
  NAND2X1 U666 ( .A(N137), .B(n404), .Y(n405) );
  NAND2X1 U667 ( .A(N136), .B(n404), .Y(n409) );
  NAND2X1 U668 ( .A(N135), .B(n404), .Y(n413) );
  NAND2X1 U669 ( .A(N134), .B(n404), .Y(n417) );
  NAND2X1 U670 ( .A(N133), .B(n404), .Y(n421) );
  NAND2X1 U671 ( .A(N132), .B(n404), .Y(n425) );
  NAND2X1 U672 ( .A(N131), .B(n404), .Y(n429) );
  NAND2X1 U673 ( .A(N138), .B(n404), .Y(n400) );
  NAND2X1 U674 ( .A(dy[7]), .B(n607), .Y(n397) );
  NAND2X1 U675 ( .A(n10), .B(n607), .Y(n360) );
  NAND2X1 U676 ( .A(N112), .B(n368), .Y(n364) );
  NAND2X1 U677 ( .A(N111), .B(n368), .Y(n369) );
  NAND2X1 U678 ( .A(N110), .B(n368), .Y(n373) );
  NAND2X1 U679 ( .A(N109), .B(n368), .Y(n377) );
  NAND2X1 U680 ( .A(N108), .B(n368), .Y(n381) );
  NAND2X1 U681 ( .A(N107), .B(n368), .Y(n385) );
  NAND2X1 U682 ( .A(N106), .B(n368), .Y(n389) );
  NAND2X1 U683 ( .A(n255), .B(n579), .Y(n363) );
  NAND2X1 U684 ( .A(N105), .B(n368), .Y(n393) );
endmodule


module screen_buffer ( clk, strb_screen, screen_cor, X0, X1, Y0, Y1 );
  input [7:0] screen_cor;
  output [7:0] X0;
  output [7:0] X1;
  output [7:0] Y0;
  output [7:0] Y1;
  input clk, strb_screen;
  wire   n3, n8, n13, n18, n23, n28, n33, n38, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n1, n2,
         n4, n5, n6, n7, n9, n10, n11, n12, n14, n15, n16, n17, n19, n20, n21,
         n22, n24, n25, n26, n27, n29, n30, n31, n32, n34, n35, n36, n37, n39,
         n40, n41, n74, n75;

  DFFPOSX1 \reg1_reg[7]  ( .D(n73), .CLK(clk), .Q(Y1[7]) );
  DFFPOSX1 \reg1_reg[15]  ( .D(n72), .CLK(clk), .Q(Y0[7]) );
  DFFPOSX1 \reg1_reg[23]  ( .D(n71), .CLK(clk), .Q(X1[7]) );
  DFFPOSX1 \reg1_reg[31]  ( .D(n70), .CLK(clk), .Q(X0[7]) );
  DFFPOSX1 \reg1_reg[6]  ( .D(n69), .CLK(clk), .Q(Y1[6]) );
  DFFPOSX1 \reg1_reg[14]  ( .D(n68), .CLK(clk), .Q(Y0[6]) );
  DFFPOSX1 \reg1_reg[22]  ( .D(n67), .CLK(clk), .Q(X1[6]) );
  DFFPOSX1 \reg1_reg[30]  ( .D(n66), .CLK(clk), .Q(X0[6]) );
  DFFPOSX1 \reg1_reg[5]  ( .D(n65), .CLK(clk), .Q(Y1[5]) );
  DFFPOSX1 \reg1_reg[13]  ( .D(n64), .CLK(clk), .Q(Y0[5]) );
  DFFPOSX1 \reg1_reg[21]  ( .D(n63), .CLK(clk), .Q(X1[5]) );
  DFFPOSX1 \reg1_reg[29]  ( .D(n62), .CLK(clk), .Q(X0[5]) );
  DFFPOSX1 \reg1_reg[4]  ( .D(n61), .CLK(clk), .Q(Y1[4]) );
  DFFPOSX1 \reg1_reg[12]  ( .D(n60), .CLK(clk), .Q(Y0[4]) );
  DFFPOSX1 \reg1_reg[20]  ( .D(n59), .CLK(clk), .Q(X1[4]) );
  DFFPOSX1 \reg1_reg[28]  ( .D(n58), .CLK(clk), .Q(X0[4]) );
  DFFPOSX1 \reg1_reg[3]  ( .D(n57), .CLK(clk), .Q(Y1[3]) );
  DFFPOSX1 \reg1_reg[11]  ( .D(n56), .CLK(clk), .Q(Y0[3]) );
  DFFPOSX1 \reg1_reg[19]  ( .D(n55), .CLK(clk), .Q(X1[3]) );
  DFFPOSX1 \reg1_reg[27]  ( .D(n54), .CLK(clk), .Q(X0[3]) );
  DFFPOSX1 \reg1_reg[2]  ( .D(n53), .CLK(clk), .Q(Y1[2]) );
  DFFPOSX1 \reg1_reg[10]  ( .D(n52), .CLK(clk), .Q(Y0[2]) );
  DFFPOSX1 \reg1_reg[18]  ( .D(n51), .CLK(clk), .Q(X1[2]) );
  DFFPOSX1 \reg1_reg[26]  ( .D(n50), .CLK(clk), .Q(X0[2]) );
  DFFPOSX1 \reg1_reg[1]  ( .D(n49), .CLK(clk), .Q(Y1[1]) );
  DFFPOSX1 \reg1_reg[9]  ( .D(n48), .CLK(clk), .Q(Y0[1]) );
  DFFPOSX1 \reg1_reg[17]  ( .D(n47), .CLK(clk), .Q(X1[1]) );
  DFFPOSX1 \reg1_reg[25]  ( .D(n46), .CLK(clk), .Q(X0[1]) );
  DFFPOSX1 \reg1_reg[0]  ( .D(n45), .CLK(clk), .Q(Y1[0]) );
  DFFPOSX1 \reg1_reg[8]  ( .D(n44), .CLK(clk), .Q(Y0[0]) );
  DFFPOSX1 \reg1_reg[16]  ( .D(n43), .CLK(clk), .Q(X1[0]) );
  DFFPOSX1 \reg1_reg[24]  ( .D(n42), .CLK(clk), .Q(X0[0]) );
  OAI21X1 U2 ( .A(n75), .B(n1), .C(n3), .Y(n42) );
  NAND2X1 U3 ( .A(X0[0]), .B(n1), .Y(n3) );
  OAI22X1 U4 ( .A(n1), .B(n74), .C(n2), .D(n75), .Y(n43) );
  OAI22X1 U6 ( .A(n1), .B(n41), .C(n2), .D(n74), .Y(n44) );
  OAI21X1 U11 ( .A(n1), .B(n40), .C(n8), .Y(n46) );
  NAND2X1 U12 ( .A(X0[1]), .B(n1), .Y(n8) );
  OAI22X1 U13 ( .A(n1), .B(n39), .C(n2), .D(n40), .Y(n47) );
  OAI22X1 U15 ( .A(n1), .B(n37), .C(n2), .D(n39), .Y(n48) );
  OAI21X1 U20 ( .A(n1), .B(n36), .C(n13), .Y(n50) );
  NAND2X1 U21 ( .A(X0[2]), .B(n1), .Y(n13) );
  OAI22X1 U22 ( .A(n1), .B(n35), .C(n2), .D(n36), .Y(n51) );
  OAI22X1 U24 ( .A(n1), .B(n34), .C(n2), .D(n35), .Y(n52) );
  OAI21X1 U29 ( .A(n1), .B(n32), .C(n18), .Y(n54) );
  NAND2X1 U30 ( .A(X0[3]), .B(n1), .Y(n18) );
  OAI22X1 U31 ( .A(n1), .B(n31), .C(n2), .D(n32), .Y(n55) );
  OAI22X1 U33 ( .A(n1), .B(n30), .C(n2), .D(n31), .Y(n56) );
  OAI21X1 U38 ( .A(n1), .B(n29), .C(n23), .Y(n58) );
  NAND2X1 U39 ( .A(X0[4]), .B(n1), .Y(n23) );
  OAI22X1 U40 ( .A(n1), .B(n27), .C(n4), .D(n29), .Y(n59) );
  OAI22X1 U42 ( .A(n1), .B(n26), .C(n4), .D(n27), .Y(n60) );
  OAI21X1 U47 ( .A(n1), .B(n25), .C(n28), .Y(n62) );
  NAND2X1 U48 ( .A(X0[5]), .B(n1), .Y(n28) );
  OAI22X1 U49 ( .A(n1), .B(n24), .C(n4), .D(n25), .Y(n63) );
  OAI22X1 U51 ( .A(n1), .B(n22), .C(n4), .D(n24), .Y(n64) );
  OAI21X1 U56 ( .A(n1), .B(n21), .C(n33), .Y(n66) );
  NAND2X1 U57 ( .A(X0[6]), .B(n1), .Y(n33) );
  OAI22X1 U58 ( .A(n1), .B(n20), .C(n4), .D(n21), .Y(n67) );
  OAI22X1 U60 ( .A(n1), .B(n19), .C(n4), .D(n20), .Y(n68) );
  OAI21X1 U65 ( .A(n1), .B(n17), .C(n38), .Y(n70) );
  NAND2X1 U66 ( .A(X0[7]), .B(n1), .Y(n38) );
  OAI22X1 U67 ( .A(n1), .B(n16), .C(n4), .D(n17), .Y(n71) );
  OAI22X1 U69 ( .A(n1), .B(n15), .C(n2), .D(n16), .Y(n72) );
  INVX4 U5 ( .A(strb_screen), .Y(n1) );
  MUX2X1 U7 ( .B(n14), .A(n15), .S(n1), .Y(n73) );
  BUFX2 U8 ( .A(strb_screen), .Y(n2) );
  BUFX2 U9 ( .A(strb_screen), .Y(n4) );
  INVX2 U10 ( .A(Y1[7]), .Y(n15) );
  INVX2 U14 ( .A(Y1[6]), .Y(n19) );
  INVX2 U16 ( .A(Y1[5]), .Y(n22) );
  INVX2 U17 ( .A(Y1[4]), .Y(n26) );
  INVX2 U18 ( .A(Y1[3]), .Y(n30) );
  INVX2 U19 ( .A(Y1[2]), .Y(n34) );
  INVX2 U23 ( .A(Y1[1]), .Y(n37) );
  INVX2 U25 ( .A(Y1[0]), .Y(n41) );
  INVX2 U26 ( .A(screen_cor[0]), .Y(n5) );
  MUX2X1 U27 ( .B(n41), .A(n5), .S(n4), .Y(n45) );
  INVX2 U28 ( .A(screen_cor[1]), .Y(n6) );
  MUX2X1 U32 ( .B(n37), .A(n6), .S(n2), .Y(n49) );
  INVX2 U34 ( .A(screen_cor[2]), .Y(n7) );
  MUX2X1 U35 ( .B(n34), .A(n7), .S(n4), .Y(n53) );
  INVX2 U36 ( .A(screen_cor[3]), .Y(n9) );
  MUX2X1 U37 ( .B(n30), .A(n9), .S(n4), .Y(n57) );
  INVX2 U41 ( .A(screen_cor[4]), .Y(n10) );
  MUX2X1 U43 ( .B(n26), .A(n10), .S(n4), .Y(n61) );
  INVX2 U44 ( .A(screen_cor[5]), .Y(n11) );
  MUX2X1 U45 ( .B(n22), .A(n11), .S(n2), .Y(n65) );
  INVX2 U46 ( .A(screen_cor[6]), .Y(n12) );
  MUX2X1 U50 ( .B(n19), .A(n12), .S(n2), .Y(n69) );
  INVX2 U52 ( .A(screen_cor[7]), .Y(n14) );
  INVX2 U53 ( .A(Y0[7]), .Y(n16) );
  INVX2 U54 ( .A(X1[7]), .Y(n17) );
  INVX2 U55 ( .A(Y0[6]), .Y(n20) );
  INVX2 U59 ( .A(X1[6]), .Y(n21) );
  INVX2 U61 ( .A(Y0[5]), .Y(n24) );
  INVX2 U62 ( .A(X1[5]), .Y(n25) );
  INVX2 U63 ( .A(Y0[4]), .Y(n27) );
  INVX2 U64 ( .A(X1[4]), .Y(n29) );
  INVX2 U68 ( .A(Y0[3]), .Y(n31) );
  INVX2 U70 ( .A(X1[3]), .Y(n32) );
  INVX2 U71 ( .A(Y0[2]), .Y(n35) );
  INVX2 U72 ( .A(X1[2]), .Y(n36) );
  INVX2 U73 ( .A(Y0[1]), .Y(n39) );
  INVX2 U74 ( .A(X1[1]), .Y(n40) );
  INVX2 U75 ( .A(Y0[0]), .Y(n74) );
  INVX2 U76 ( .A(X1[0]), .Y(n75) );
endmodule


module world_matrix_buffer ( strb_matrix, databus_out, clk, row_sel, row );
  input [15:0] databus_out;
  input [1:0] row_sel;
  output [63:0] row;
  input strb_matrix, clk;
  wire   n134, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n406, n420, n421, n422, n436, n437, n438, n452,
         n453, n454, n468, n469, n470, n484, n485, n486, n500, n501, n502,
         n516, n517, n518, n532, n533, n534, n548, n549, n550, n564, n565,
         n566, n580, n581, n582, n596, n597, n598, n612, n613, n614, n628,
         n629, n630, n644, n645, n646, n660, n661, n662, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n135, n148, n149,
         n150, n165, n166, n167, n182, n183, n184, n199, n200, n201, n216,
         n217, n218, n233, n234, n235, n250, n251, n252, n267, n268, n269,
         n284, n285, n286, n301, n302, n303, n318, n319, n320, n335, n336,
         n337, n352, n353, n354, n369, n370, n371, n386, n387, n388, n403,
         n404, n405, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804;
  wire   [255:0] regg;
  tri   [15:0] databus_out;

  DFFPOSX1 \regg_reg[15]  ( .D(n662), .CLK(clk), .Q(regg[15]) );
  DFFPOSX1 \regg_reg[31]  ( .D(n661), .CLK(clk), .Q(regg[31]) );
  DFFPOSX1 \regg_reg[47]  ( .D(n660), .CLK(clk), .Q(regg[47]) );
  DFFPOSX1 \regg_reg[63]  ( .D(n756), .CLK(clk), .Q(regg[63]) );
  DFFPOSX1 \regg_reg[79]  ( .D(n755), .CLK(clk), .Q(regg[79]) );
  DFFPOSX1 \regg_reg[95]  ( .D(n754), .CLK(clk), .Q(regg[95]) );
  DFFPOSX1 \regg_reg[111]  ( .D(n753), .CLK(clk), .Q(regg[111]) );
  DFFPOSX1 \regg_reg[127]  ( .D(n752), .CLK(clk), .Q(regg[127]) );
  DFFPOSX1 \regg_reg[143]  ( .D(n751), .CLK(clk), .Q(regg[143]) );
  DFFPOSX1 \regg_reg[159]  ( .D(n750), .CLK(clk), .Q(regg[159]) );
  DFFPOSX1 \regg_reg[175]  ( .D(n749), .CLK(clk), .Q(regg[175]) );
  DFFPOSX1 \regg_reg[191]  ( .D(n748), .CLK(clk), .Q(regg[191]) );
  DFFPOSX1 \regg_reg[207]  ( .D(n747), .CLK(clk), .Q(regg[207]) );
  DFFPOSX1 \regg_reg[223]  ( .D(n746), .CLK(clk), .Q(regg[223]) );
  DFFPOSX1 \regg_reg[239]  ( .D(n745), .CLK(clk), .Q(regg[239]) );
  DFFPOSX1 \regg_reg[255]  ( .D(n744), .CLK(clk), .Q(regg[255]) );
  DFFPOSX1 \regg_reg[14]  ( .D(n646), .CLK(clk), .Q(regg[14]) );
  DFFPOSX1 \regg_reg[30]  ( .D(n645), .CLK(clk), .Q(regg[30]) );
  DFFPOSX1 \regg_reg[46]  ( .D(n644), .CLK(clk), .Q(regg[46]) );
  DFFPOSX1 \regg_reg[62]  ( .D(n743), .CLK(clk), .Q(regg[62]) );
  DFFPOSX1 \regg_reg[78]  ( .D(n742), .CLK(clk), .Q(regg[78]) );
  DFFPOSX1 \regg_reg[94]  ( .D(n741), .CLK(clk), .Q(regg[94]) );
  DFFPOSX1 \regg_reg[110]  ( .D(n740), .CLK(clk), .Q(regg[110]) );
  DFFPOSX1 \regg_reg[126]  ( .D(n739), .CLK(clk), .Q(regg[126]) );
  DFFPOSX1 \regg_reg[142]  ( .D(n738), .CLK(clk), .Q(regg[142]) );
  DFFPOSX1 \regg_reg[158]  ( .D(n737), .CLK(clk), .Q(regg[158]) );
  DFFPOSX1 \regg_reg[174]  ( .D(n736), .CLK(clk), .Q(regg[174]) );
  DFFPOSX1 \regg_reg[190]  ( .D(n735), .CLK(clk), .Q(regg[190]) );
  DFFPOSX1 \regg_reg[206]  ( .D(n734), .CLK(clk), .Q(regg[206]) );
  DFFPOSX1 \regg_reg[222]  ( .D(n733), .CLK(clk), .Q(regg[222]) );
  DFFPOSX1 \regg_reg[238]  ( .D(n732), .CLK(clk), .Q(regg[238]) );
  DFFPOSX1 \regg_reg[254]  ( .D(n731), .CLK(clk), .Q(regg[254]) );
  DFFPOSX1 \regg_reg[13]  ( .D(n630), .CLK(clk), .Q(regg[13]) );
  DFFPOSX1 \regg_reg[29]  ( .D(n629), .CLK(clk), .Q(regg[29]) );
  DFFPOSX1 \regg_reg[45]  ( .D(n628), .CLK(clk), .Q(regg[45]) );
  DFFPOSX1 \regg_reg[61]  ( .D(n730), .CLK(clk), .Q(regg[61]) );
  DFFPOSX1 \regg_reg[77]  ( .D(n729), .CLK(clk), .Q(regg[77]) );
  DFFPOSX1 \regg_reg[93]  ( .D(n728), .CLK(clk), .Q(regg[93]) );
  DFFPOSX1 \regg_reg[109]  ( .D(n727), .CLK(clk), .Q(regg[109]) );
  DFFPOSX1 \regg_reg[125]  ( .D(n726), .CLK(clk), .Q(regg[125]) );
  DFFPOSX1 \regg_reg[141]  ( .D(n725), .CLK(clk), .Q(regg[141]) );
  DFFPOSX1 \regg_reg[157]  ( .D(n724), .CLK(clk), .Q(regg[157]) );
  DFFPOSX1 \regg_reg[173]  ( .D(n723), .CLK(clk), .Q(regg[173]) );
  DFFPOSX1 \regg_reg[189]  ( .D(n722), .CLK(clk), .Q(regg[189]) );
  DFFPOSX1 \regg_reg[205]  ( .D(n721), .CLK(clk), .Q(regg[205]) );
  DFFPOSX1 \regg_reg[221]  ( .D(n720), .CLK(clk), .Q(regg[221]) );
  DFFPOSX1 \regg_reg[237]  ( .D(n719), .CLK(clk), .Q(regg[237]) );
  DFFPOSX1 \regg_reg[253]  ( .D(n718), .CLK(clk), .Q(regg[253]) );
  DFFPOSX1 \regg_reg[12]  ( .D(n614), .CLK(clk), .Q(regg[12]) );
  DFFPOSX1 \regg_reg[28]  ( .D(n613), .CLK(clk), .Q(regg[28]) );
  DFFPOSX1 \regg_reg[44]  ( .D(n612), .CLK(clk), .Q(regg[44]) );
  DFFPOSX1 \regg_reg[60]  ( .D(n717), .CLK(clk), .Q(regg[60]) );
  DFFPOSX1 \regg_reg[76]  ( .D(n716), .CLK(clk), .Q(regg[76]) );
  DFFPOSX1 \regg_reg[92]  ( .D(n715), .CLK(clk), .Q(regg[92]) );
  DFFPOSX1 \regg_reg[108]  ( .D(n714), .CLK(clk), .Q(regg[108]) );
  DFFPOSX1 \regg_reg[124]  ( .D(n713), .CLK(clk), .Q(regg[124]) );
  DFFPOSX1 \regg_reg[140]  ( .D(n712), .CLK(clk), .Q(regg[140]) );
  DFFPOSX1 \regg_reg[156]  ( .D(n711), .CLK(clk), .Q(regg[156]) );
  DFFPOSX1 \regg_reg[172]  ( .D(n710), .CLK(clk), .Q(regg[172]) );
  DFFPOSX1 \regg_reg[188]  ( .D(n709), .CLK(clk), .Q(regg[188]) );
  DFFPOSX1 \regg_reg[204]  ( .D(n708), .CLK(clk), .Q(regg[204]) );
  DFFPOSX1 \regg_reg[220]  ( .D(n707), .CLK(clk), .Q(regg[220]) );
  DFFPOSX1 \regg_reg[236]  ( .D(n706), .CLK(clk), .Q(regg[236]) );
  DFFPOSX1 \regg_reg[252]  ( .D(n705), .CLK(clk), .Q(regg[252]) );
  DFFPOSX1 \regg_reg[11]  ( .D(n598), .CLK(clk), .Q(regg[11]) );
  DFFPOSX1 \regg_reg[27]  ( .D(n597), .CLK(clk), .Q(regg[27]) );
  DFFPOSX1 \regg_reg[43]  ( .D(n596), .CLK(clk), .Q(regg[43]) );
  DFFPOSX1 \regg_reg[59]  ( .D(n704), .CLK(clk), .Q(regg[59]) );
  DFFPOSX1 \regg_reg[75]  ( .D(n703), .CLK(clk), .Q(regg[75]) );
  DFFPOSX1 \regg_reg[91]  ( .D(n702), .CLK(clk), .Q(regg[91]) );
  DFFPOSX1 \regg_reg[107]  ( .D(n701), .CLK(clk), .Q(regg[107]) );
  DFFPOSX1 \regg_reg[123]  ( .D(n700), .CLK(clk), .Q(regg[123]) );
  DFFPOSX1 \regg_reg[139]  ( .D(n699), .CLK(clk), .Q(regg[139]) );
  DFFPOSX1 \regg_reg[155]  ( .D(n698), .CLK(clk), .Q(regg[155]) );
  DFFPOSX1 \regg_reg[171]  ( .D(n697), .CLK(clk), .Q(regg[171]) );
  DFFPOSX1 \regg_reg[187]  ( .D(n696), .CLK(clk), .Q(regg[187]) );
  DFFPOSX1 \regg_reg[203]  ( .D(n695), .CLK(clk), .Q(regg[203]) );
  DFFPOSX1 \regg_reg[219]  ( .D(n694), .CLK(clk), .Q(regg[219]) );
  DFFPOSX1 \regg_reg[235]  ( .D(n693), .CLK(clk), .Q(regg[235]) );
  DFFPOSX1 \regg_reg[251]  ( .D(n692), .CLK(clk), .Q(regg[251]) );
  DFFPOSX1 \regg_reg[10]  ( .D(n582), .CLK(clk), .Q(regg[10]) );
  DFFPOSX1 \regg_reg[26]  ( .D(n581), .CLK(clk), .Q(regg[26]) );
  DFFPOSX1 \regg_reg[42]  ( .D(n580), .CLK(clk), .Q(regg[42]) );
  DFFPOSX1 \regg_reg[58]  ( .D(n691), .CLK(clk), .Q(regg[58]) );
  DFFPOSX1 \regg_reg[74]  ( .D(n690), .CLK(clk), .Q(regg[74]) );
  DFFPOSX1 \regg_reg[90]  ( .D(n689), .CLK(clk), .Q(regg[90]) );
  DFFPOSX1 \regg_reg[106]  ( .D(n688), .CLK(clk), .Q(regg[106]) );
  DFFPOSX1 \regg_reg[122]  ( .D(n687), .CLK(clk), .Q(regg[122]) );
  DFFPOSX1 \regg_reg[138]  ( .D(n686), .CLK(clk), .Q(regg[138]) );
  DFFPOSX1 \regg_reg[154]  ( .D(n685), .CLK(clk), .Q(regg[154]) );
  DFFPOSX1 \regg_reg[170]  ( .D(n684), .CLK(clk), .Q(regg[170]) );
  DFFPOSX1 \regg_reg[186]  ( .D(n683), .CLK(clk), .Q(regg[186]) );
  DFFPOSX1 \regg_reg[202]  ( .D(n682), .CLK(clk), .Q(regg[202]) );
  DFFPOSX1 \regg_reg[218]  ( .D(n681), .CLK(clk), .Q(regg[218]) );
  DFFPOSX1 \regg_reg[234]  ( .D(n680), .CLK(clk), .Q(regg[234]) );
  DFFPOSX1 \regg_reg[250]  ( .D(n679), .CLK(clk), .Q(regg[250]) );
  DFFPOSX1 \regg_reg[9]  ( .D(n566), .CLK(clk), .Q(regg[9]) );
  DFFPOSX1 \regg_reg[25]  ( .D(n565), .CLK(clk), .Q(regg[25]) );
  DFFPOSX1 \regg_reg[41]  ( .D(n564), .CLK(clk), .Q(regg[41]) );
  DFFPOSX1 \regg_reg[57]  ( .D(n678), .CLK(clk), .Q(regg[57]) );
  DFFPOSX1 \regg_reg[73]  ( .D(n677), .CLK(clk), .Q(regg[73]) );
  DFFPOSX1 \regg_reg[89]  ( .D(n676), .CLK(clk), .Q(regg[89]) );
  DFFPOSX1 \regg_reg[105]  ( .D(n675), .CLK(clk), .Q(regg[105]) );
  DFFPOSX1 \regg_reg[121]  ( .D(n674), .CLK(clk), .Q(regg[121]) );
  DFFPOSX1 \regg_reg[137]  ( .D(n673), .CLK(clk), .Q(regg[137]) );
  DFFPOSX1 \regg_reg[153]  ( .D(n672), .CLK(clk), .Q(regg[153]) );
  DFFPOSX1 \regg_reg[169]  ( .D(n671), .CLK(clk), .Q(regg[169]) );
  DFFPOSX1 \regg_reg[185]  ( .D(n670), .CLK(clk), .Q(regg[185]) );
  DFFPOSX1 \regg_reg[201]  ( .D(n669), .CLK(clk), .Q(regg[201]) );
  DFFPOSX1 \regg_reg[217]  ( .D(n668), .CLK(clk), .Q(regg[217]) );
  DFFPOSX1 \regg_reg[233]  ( .D(n667), .CLK(clk), .Q(regg[233]) );
  DFFPOSX1 \regg_reg[249]  ( .D(n666), .CLK(clk), .Q(regg[249]) );
  DFFPOSX1 \regg_reg[8]  ( .D(n550), .CLK(clk), .Q(regg[8]) );
  DFFPOSX1 \regg_reg[24]  ( .D(n549), .CLK(clk), .Q(regg[24]) );
  DFFPOSX1 \regg_reg[40]  ( .D(n548), .CLK(clk), .Q(regg[40]) );
  DFFPOSX1 \regg_reg[56]  ( .D(n665), .CLK(clk), .Q(regg[56]) );
  DFFPOSX1 \regg_reg[72]  ( .D(n664), .CLK(clk), .Q(regg[72]) );
  DFFPOSX1 \regg_reg[88]  ( .D(n663), .CLK(clk), .Q(regg[88]) );
  DFFPOSX1 \regg_reg[104]  ( .D(n659), .CLK(clk), .Q(regg[104]) );
  DFFPOSX1 \regg_reg[120]  ( .D(n658), .CLK(clk), .Q(regg[120]) );
  DFFPOSX1 \regg_reg[136]  ( .D(n657), .CLK(clk), .Q(regg[136]) );
  DFFPOSX1 \regg_reg[152]  ( .D(n656), .CLK(clk), .Q(regg[152]) );
  DFFPOSX1 \regg_reg[168]  ( .D(n655), .CLK(clk), .Q(regg[168]) );
  DFFPOSX1 \regg_reg[184]  ( .D(n654), .CLK(clk), .Q(regg[184]) );
  DFFPOSX1 \regg_reg[200]  ( .D(n653), .CLK(clk), .Q(regg[200]) );
  DFFPOSX1 \regg_reg[216]  ( .D(n652), .CLK(clk), .Q(regg[216]) );
  DFFPOSX1 \regg_reg[232]  ( .D(n651), .CLK(clk), .Q(regg[232]) );
  DFFPOSX1 \regg_reg[248]  ( .D(n650), .CLK(clk), .Q(regg[248]) );
  DFFPOSX1 \regg_reg[7]  ( .D(n534), .CLK(clk), .Q(regg[7]) );
  DFFPOSX1 \regg_reg[23]  ( .D(n533), .CLK(clk), .Q(regg[23]) );
  DFFPOSX1 \regg_reg[39]  ( .D(n532), .CLK(clk), .Q(regg[39]) );
  DFFPOSX1 \regg_reg[55]  ( .D(n649), .CLK(clk), .Q(regg[55]) );
  DFFPOSX1 \regg_reg[71]  ( .D(n648), .CLK(clk), .Q(regg[71]) );
  DFFPOSX1 \regg_reg[87]  ( .D(n647), .CLK(clk), .Q(regg[87]) );
  DFFPOSX1 \regg_reg[103]  ( .D(n643), .CLK(clk), .Q(regg[103]) );
  DFFPOSX1 \regg_reg[119]  ( .D(n642), .CLK(clk), .Q(regg[119]) );
  DFFPOSX1 \regg_reg[135]  ( .D(n641), .CLK(clk), .Q(regg[135]) );
  DFFPOSX1 \regg_reg[151]  ( .D(n640), .CLK(clk), .Q(regg[151]) );
  DFFPOSX1 \regg_reg[167]  ( .D(n639), .CLK(clk), .Q(regg[167]) );
  DFFPOSX1 \regg_reg[183]  ( .D(n638), .CLK(clk), .Q(regg[183]) );
  DFFPOSX1 \regg_reg[199]  ( .D(n637), .CLK(clk), .Q(regg[199]) );
  DFFPOSX1 \regg_reg[215]  ( .D(n636), .CLK(clk), .Q(regg[215]) );
  DFFPOSX1 \regg_reg[231]  ( .D(n635), .CLK(clk), .Q(regg[231]) );
  DFFPOSX1 \regg_reg[247]  ( .D(n634), .CLK(clk), .Q(regg[247]) );
  DFFPOSX1 \regg_reg[6]  ( .D(n518), .CLK(clk), .Q(regg[6]) );
  DFFPOSX1 \regg_reg[22]  ( .D(n517), .CLK(clk), .Q(regg[22]) );
  DFFPOSX1 \regg_reg[38]  ( .D(n516), .CLK(clk), .Q(regg[38]) );
  DFFPOSX1 \regg_reg[54]  ( .D(n633), .CLK(clk), .Q(regg[54]) );
  DFFPOSX1 \regg_reg[70]  ( .D(n632), .CLK(clk), .Q(regg[70]) );
  DFFPOSX1 \regg_reg[86]  ( .D(n631), .CLK(clk), .Q(regg[86]) );
  DFFPOSX1 \regg_reg[102]  ( .D(n627), .CLK(clk), .Q(regg[102]) );
  DFFPOSX1 \regg_reg[118]  ( .D(n626), .CLK(clk), .Q(regg[118]) );
  DFFPOSX1 \regg_reg[134]  ( .D(n625), .CLK(clk), .Q(regg[134]) );
  DFFPOSX1 \regg_reg[150]  ( .D(n624), .CLK(clk), .Q(regg[150]) );
  DFFPOSX1 \regg_reg[166]  ( .D(n623), .CLK(clk), .Q(regg[166]) );
  DFFPOSX1 \regg_reg[182]  ( .D(n622), .CLK(clk), .Q(regg[182]) );
  DFFPOSX1 \regg_reg[198]  ( .D(n621), .CLK(clk), .Q(regg[198]) );
  DFFPOSX1 \regg_reg[214]  ( .D(n620), .CLK(clk), .Q(regg[214]) );
  DFFPOSX1 \regg_reg[230]  ( .D(n619), .CLK(clk), .Q(regg[230]) );
  DFFPOSX1 \regg_reg[246]  ( .D(n618), .CLK(clk), .Q(regg[246]) );
  DFFPOSX1 \regg_reg[5]  ( .D(n502), .CLK(clk), .Q(regg[5]) );
  DFFPOSX1 \regg_reg[21]  ( .D(n501), .CLK(clk), .Q(regg[21]) );
  DFFPOSX1 \regg_reg[37]  ( .D(n500), .CLK(clk), .Q(regg[37]) );
  DFFPOSX1 \regg_reg[53]  ( .D(n617), .CLK(clk), .Q(regg[53]) );
  DFFPOSX1 \regg_reg[69]  ( .D(n616), .CLK(clk), .Q(regg[69]) );
  DFFPOSX1 \regg_reg[85]  ( .D(n615), .CLK(clk), .Q(regg[85]) );
  DFFPOSX1 \regg_reg[101]  ( .D(n611), .CLK(clk), .Q(regg[101]) );
  DFFPOSX1 \regg_reg[117]  ( .D(n610), .CLK(clk), .Q(regg[117]) );
  DFFPOSX1 \regg_reg[133]  ( .D(n609), .CLK(clk), .Q(regg[133]) );
  DFFPOSX1 \regg_reg[149]  ( .D(n608), .CLK(clk), .Q(regg[149]) );
  DFFPOSX1 \regg_reg[165]  ( .D(n607), .CLK(clk), .Q(regg[165]) );
  DFFPOSX1 \regg_reg[181]  ( .D(n606), .CLK(clk), .Q(regg[181]) );
  DFFPOSX1 \regg_reg[197]  ( .D(n605), .CLK(clk), .Q(regg[197]) );
  DFFPOSX1 \regg_reg[213]  ( .D(n604), .CLK(clk), .Q(regg[213]) );
  DFFPOSX1 \regg_reg[229]  ( .D(n603), .CLK(clk), .Q(regg[229]) );
  DFFPOSX1 \regg_reg[245]  ( .D(n602), .CLK(clk), .Q(regg[245]) );
  DFFPOSX1 \regg_reg[4]  ( .D(n486), .CLK(clk), .Q(regg[4]) );
  DFFPOSX1 \regg_reg[20]  ( .D(n485), .CLK(clk), .Q(regg[20]) );
  DFFPOSX1 \regg_reg[36]  ( .D(n484), .CLK(clk), .Q(regg[36]) );
  DFFPOSX1 \regg_reg[52]  ( .D(n601), .CLK(clk), .Q(regg[52]) );
  DFFPOSX1 \regg_reg[68]  ( .D(n600), .CLK(clk), .Q(regg[68]) );
  DFFPOSX1 \regg_reg[84]  ( .D(n599), .CLK(clk), .Q(regg[84]) );
  DFFPOSX1 \regg_reg[100]  ( .D(n595), .CLK(clk), .Q(regg[100]) );
  DFFPOSX1 \regg_reg[116]  ( .D(n594), .CLK(clk), .Q(regg[116]) );
  DFFPOSX1 \regg_reg[132]  ( .D(n593), .CLK(clk), .Q(regg[132]) );
  DFFPOSX1 \regg_reg[148]  ( .D(n592), .CLK(clk), .Q(regg[148]) );
  DFFPOSX1 \regg_reg[164]  ( .D(n591), .CLK(clk), .Q(regg[164]) );
  DFFPOSX1 \regg_reg[180]  ( .D(n590), .CLK(clk), .Q(regg[180]) );
  DFFPOSX1 \regg_reg[196]  ( .D(n589), .CLK(clk), .Q(regg[196]) );
  DFFPOSX1 \regg_reg[212]  ( .D(n588), .CLK(clk), .Q(regg[212]) );
  DFFPOSX1 \regg_reg[228]  ( .D(n587), .CLK(clk), .Q(regg[228]) );
  DFFPOSX1 \regg_reg[244]  ( .D(n586), .CLK(clk), .Q(regg[244]) );
  DFFPOSX1 \regg_reg[3]  ( .D(n470), .CLK(clk), .Q(regg[3]) );
  DFFPOSX1 \regg_reg[19]  ( .D(n469), .CLK(clk), .Q(regg[19]) );
  DFFPOSX1 \regg_reg[35]  ( .D(n468), .CLK(clk), .Q(regg[35]) );
  DFFPOSX1 \regg_reg[51]  ( .D(n585), .CLK(clk), .Q(regg[51]) );
  DFFPOSX1 \regg_reg[67]  ( .D(n584), .CLK(clk), .Q(regg[67]) );
  DFFPOSX1 \regg_reg[83]  ( .D(n583), .CLK(clk), .Q(regg[83]) );
  DFFPOSX1 \regg_reg[99]  ( .D(n579), .CLK(clk), .Q(regg[99]) );
  DFFPOSX1 \regg_reg[115]  ( .D(n578), .CLK(clk), .Q(regg[115]) );
  DFFPOSX1 \regg_reg[131]  ( .D(n577), .CLK(clk), .Q(regg[131]) );
  DFFPOSX1 \regg_reg[147]  ( .D(n576), .CLK(clk), .Q(regg[147]) );
  DFFPOSX1 \regg_reg[163]  ( .D(n575), .CLK(clk), .Q(regg[163]) );
  DFFPOSX1 \regg_reg[179]  ( .D(n574), .CLK(clk), .Q(regg[179]) );
  DFFPOSX1 \regg_reg[195]  ( .D(n573), .CLK(clk), .Q(regg[195]) );
  DFFPOSX1 \regg_reg[211]  ( .D(n572), .CLK(clk), .Q(regg[211]) );
  DFFPOSX1 \regg_reg[227]  ( .D(n571), .CLK(clk), .Q(regg[227]) );
  DFFPOSX1 \regg_reg[243]  ( .D(n570), .CLK(clk), .Q(regg[243]) );
  DFFPOSX1 \regg_reg[2]  ( .D(n454), .CLK(clk), .Q(regg[2]) );
  DFFPOSX1 \regg_reg[18]  ( .D(n453), .CLK(clk), .Q(regg[18]) );
  DFFPOSX1 \regg_reg[34]  ( .D(n452), .CLK(clk), .Q(regg[34]) );
  DFFPOSX1 \regg_reg[50]  ( .D(n569), .CLK(clk), .Q(regg[50]) );
  DFFPOSX1 \regg_reg[66]  ( .D(n568), .CLK(clk), .Q(regg[66]) );
  DFFPOSX1 \regg_reg[82]  ( .D(n567), .CLK(clk), .Q(regg[82]) );
  DFFPOSX1 \regg_reg[98]  ( .D(n563), .CLK(clk), .Q(regg[98]) );
  DFFPOSX1 \regg_reg[114]  ( .D(n562), .CLK(clk), .Q(regg[114]) );
  DFFPOSX1 \regg_reg[130]  ( .D(n561), .CLK(clk), .Q(regg[130]) );
  DFFPOSX1 \regg_reg[146]  ( .D(n560), .CLK(clk), .Q(regg[146]) );
  DFFPOSX1 \regg_reg[162]  ( .D(n559), .CLK(clk), .Q(regg[162]) );
  DFFPOSX1 \regg_reg[178]  ( .D(n558), .CLK(clk), .Q(regg[178]) );
  DFFPOSX1 \regg_reg[194]  ( .D(n557), .CLK(clk), .Q(regg[194]) );
  DFFPOSX1 \regg_reg[210]  ( .D(n556), .CLK(clk), .Q(regg[210]) );
  DFFPOSX1 \regg_reg[226]  ( .D(n555), .CLK(clk), .Q(regg[226]) );
  DFFPOSX1 \regg_reg[242]  ( .D(n554), .CLK(clk), .Q(regg[242]) );
  DFFPOSX1 \regg_reg[1]  ( .D(n438), .CLK(clk), .Q(regg[1]) );
  DFFPOSX1 \regg_reg[17]  ( .D(n437), .CLK(clk), .Q(regg[17]) );
  DFFPOSX1 \regg_reg[33]  ( .D(n436), .CLK(clk), .Q(regg[33]) );
  DFFPOSX1 \regg_reg[49]  ( .D(n553), .CLK(clk), .Q(regg[49]) );
  DFFPOSX1 \regg_reg[65]  ( .D(n552), .CLK(clk), .Q(regg[65]) );
  DFFPOSX1 \regg_reg[81]  ( .D(n551), .CLK(clk), .Q(regg[81]) );
  DFFPOSX1 \regg_reg[97]  ( .D(n547), .CLK(clk), .Q(regg[97]) );
  DFFPOSX1 \regg_reg[113]  ( .D(n546), .CLK(clk), .Q(regg[113]) );
  DFFPOSX1 \regg_reg[129]  ( .D(n545), .CLK(clk), .Q(regg[129]) );
  DFFPOSX1 \regg_reg[145]  ( .D(n544), .CLK(clk), .Q(regg[145]) );
  DFFPOSX1 \regg_reg[161]  ( .D(n543), .CLK(clk), .Q(regg[161]) );
  DFFPOSX1 \regg_reg[177]  ( .D(n542), .CLK(clk), .Q(regg[177]) );
  DFFPOSX1 \regg_reg[193]  ( .D(n541), .CLK(clk), .Q(regg[193]) );
  DFFPOSX1 \regg_reg[209]  ( .D(n540), .CLK(clk), .Q(regg[209]) );
  DFFPOSX1 \regg_reg[225]  ( .D(n539), .CLK(clk), .Q(regg[225]) );
  DFFPOSX1 \regg_reg[241]  ( .D(n538), .CLK(clk), .Q(regg[241]) );
  DFFPOSX1 \regg_reg[0]  ( .D(n422), .CLK(clk), .Q(regg[0]) );
  DFFPOSX1 \regg_reg[16]  ( .D(n421), .CLK(clk), .Q(regg[16]) );
  DFFPOSX1 \regg_reg[32]  ( .D(n420), .CLK(clk), .Q(regg[32]) );
  DFFPOSX1 \regg_reg[48]  ( .D(n537), .CLK(clk), .Q(regg[48]) );
  DFFPOSX1 \regg_reg[64]  ( .D(n536), .CLK(clk), .Q(regg[64]) );
  DFFPOSX1 \regg_reg[80]  ( .D(n535), .CLK(clk), .Q(regg[80]) );
  DFFPOSX1 \regg_reg[96]  ( .D(n531), .CLK(clk), .Q(regg[96]) );
  DFFPOSX1 \regg_reg[112]  ( .D(n530), .CLK(clk), .Q(regg[112]) );
  DFFPOSX1 \regg_reg[128]  ( .D(n529), .CLK(clk), .Q(regg[128]) );
  DFFPOSX1 \regg_reg[144]  ( .D(n528), .CLK(clk), .Q(regg[144]) );
  DFFPOSX1 \regg_reg[160]  ( .D(n527), .CLK(clk), .Q(regg[160]) );
  DFFPOSX1 \regg_reg[176]  ( .D(n526), .CLK(clk), .Q(regg[176]) );
  DFFPOSX1 \regg_reg[192]  ( .D(n525), .CLK(clk), .Q(regg[192]) );
  DFFPOSX1 \regg_reg[208]  ( .D(n524), .CLK(clk), .Q(regg[208]) );
  DFFPOSX1 \regg_reg[224]  ( .D(n523), .CLK(clk), .Q(regg[224]) );
  DFFPOSX1 \regg_reg[240]  ( .D(n522), .CLK(clk), .Q(regg[240]) );
  AOI22X1 U200 ( .A(n96), .B(regg[240]), .C(regg[224]), .D(n46), .Y(n134) );
  AOI22X1 U202 ( .A(n96), .B(regg[224]), .C(regg[208]), .D(n46), .Y(n136) );
  AOI22X1 U204 ( .A(n96), .B(regg[208]), .C(regg[192]), .D(n46), .Y(n137) );
  AOI22X1 U206 ( .A(n95), .B(regg[192]), .C(regg[176]), .D(n46), .Y(n138) );
  AOI22X1 U208 ( .A(n95), .B(regg[176]), .C(regg[160]), .D(n47), .Y(n139) );
  AOI22X1 U210 ( .A(n94), .B(regg[160]), .C(regg[144]), .D(n47), .Y(n140) );
  AOI22X1 U212 ( .A(n94), .B(regg[144]), .C(regg[128]), .D(n47), .Y(n141) );
  AOI22X1 U214 ( .A(n92), .B(regg[128]), .C(regg[112]), .D(n47), .Y(n142) );
  AOI22X1 U216 ( .A(regg[96]), .B(n60), .C(n75), .D(regg[112]), .Y(n143) );
  AOI22X1 U218 ( .A(n92), .B(regg[96]), .C(regg[80]), .D(n47), .Y(n144) );
  AOI22X1 U220 ( .A(n92), .B(regg[80]), .C(regg[64]), .D(n47), .Y(n145) );
  AOI22X1 U222 ( .A(n91), .B(regg[64]), .C(regg[48]), .D(n46), .Y(n146) );
  AOI22X1 U224 ( .A(n91), .B(regg[48]), .C(regg[32]), .D(n46), .Y(n147) );
  OAI22X1 U225 ( .A(n62), .B(n804), .C(n803), .D(n73), .Y(n420) );
  OAI22X1 U227 ( .A(n62), .B(n803), .C(n802), .D(n71), .Y(n421) );
  OAI21X1 U229 ( .A(n65), .B(n802), .C(n151), .Y(n422) );
  NAND2X1 U230 ( .A(databus_out[0]), .B(n64), .Y(n151) );
  AOI22X1 U233 ( .A(n91), .B(regg[241]), .C(regg[225]), .D(n47), .Y(n152) );
  AOI22X1 U235 ( .A(n89), .B(regg[225]), .C(regg[209]), .D(n57), .Y(n153) );
  AOI22X1 U237 ( .A(n88), .B(regg[209]), .C(regg[193]), .D(n48), .Y(n154) );
  AOI22X1 U239 ( .A(n88), .B(regg[193]), .C(regg[177]), .D(n48), .Y(n155) );
  AOI22X1 U241 ( .A(n88), .B(regg[177]), .C(regg[161]), .D(n48), .Y(n156) );
  AOI22X1 U243 ( .A(n87), .B(regg[161]), .C(regg[145]), .D(n48), .Y(n157) );
  AOI22X1 U245 ( .A(n86), .B(regg[145]), .C(regg[129]), .D(n48), .Y(n158) );
  AOI22X1 U247 ( .A(n85), .B(regg[129]), .C(regg[113]), .D(n48), .Y(n159) );
  AOI22X1 U249 ( .A(regg[97]), .B(n60), .C(n77), .D(regg[113]), .Y(n160) );
  AOI22X1 U251 ( .A(n85), .B(regg[97]), .C(regg[81]), .D(n57), .Y(n161) );
  AOI22X1 U253 ( .A(n85), .B(regg[81]), .C(regg[65]), .D(n48), .Y(n162) );
  AOI22X1 U255 ( .A(n84), .B(regg[65]), .C(regg[49]), .D(n57), .Y(n163) );
  AOI22X1 U257 ( .A(n83), .B(regg[49]), .C(regg[33]), .D(n58), .Y(n164) );
  OAI22X1 U258 ( .A(n64), .B(n801), .C(n800), .D(n73), .Y(n436) );
  OAI22X1 U260 ( .A(n799), .B(n79), .C(n62), .D(n800), .Y(n437) );
  OAI21X1 U262 ( .A(n64), .B(n799), .C(n168), .Y(n438) );
  NAND2X1 U263 ( .A(databus_out[1]), .B(n65), .Y(n168) );
  AOI22X1 U266 ( .A(n82), .B(regg[242]), .C(regg[226]), .D(n49), .Y(n169) );
  AOI22X1 U268 ( .A(n82), .B(regg[226]), .C(regg[210]), .D(n49), .Y(n170) );
  AOI22X1 U270 ( .A(n81), .B(regg[210]), .C(regg[194]), .D(n58), .Y(n171) );
  AOI22X1 U272 ( .A(n81), .B(regg[194]), .C(regg[178]), .D(n49), .Y(n172) );
  AOI22X1 U274 ( .A(n80), .B(regg[178]), .C(regg[162]), .D(n49), .Y(n173) );
  AOI22X1 U276 ( .A(n80), .B(regg[162]), .C(regg[146]), .D(n49), .Y(n174) );
  AOI22X1 U278 ( .A(n79), .B(regg[146]), .C(regg[130]), .D(n49), .Y(n175) );
  AOI22X1 U280 ( .A(n80), .B(regg[130]), .C(regg[114]), .D(n49), .Y(n176) );
  AOI22X1 U282 ( .A(regg[98]), .B(n61), .C(n77), .D(regg[114]), .Y(n177) );
  AOI22X1 U284 ( .A(n80), .B(regg[98]), .C(regg[82]), .D(n49), .Y(n178) );
  AOI22X1 U286 ( .A(n80), .B(regg[82]), .C(regg[66]), .D(n50), .Y(n179) );
  AOI22X1 U288 ( .A(n81), .B(regg[66]), .C(regg[50]), .D(n50), .Y(n180) );
  AOI22X1 U290 ( .A(n81), .B(regg[50]), .C(regg[34]), .D(n58), .Y(n181) );
  OAI22X1 U291 ( .A(n63), .B(n798), .C(n797), .D(n74), .Y(n452) );
  OAI22X1 U293 ( .A(n796), .B(n78), .C(n62), .D(n797), .Y(n453) );
  OAI21X1 U295 ( .A(n64), .B(n796), .C(n185), .Y(n454) );
  NAND2X1 U296 ( .A(databus_out[2]), .B(n65), .Y(n185) );
  AOI22X1 U299 ( .A(n81), .B(regg[243]), .C(regg[227]), .D(n59), .Y(n186) );
  AOI22X1 U301 ( .A(n82), .B(regg[227]), .C(regg[211]), .D(n59), .Y(n187) );
  AOI22X1 U303 ( .A(n82), .B(regg[211]), .C(regg[195]), .D(n50), .Y(n188) );
  AOI22X1 U305 ( .A(n82), .B(regg[195]), .C(regg[179]), .D(n50), .Y(n189) );
  AOI22X1 U307 ( .A(n83), .B(regg[179]), .C(regg[163]), .D(n50), .Y(n190) );
  AOI22X1 U309 ( .A(n83), .B(regg[163]), .C(regg[147]), .D(n59), .Y(n191) );
  AOI22X1 U311 ( .A(n83), .B(regg[147]), .C(regg[131]), .D(n51), .Y(n192) );
  AOI22X1 U313 ( .A(n83), .B(regg[131]), .C(regg[115]), .D(n51), .Y(n193) );
  AOI22X1 U315 ( .A(regg[99]), .B(n61), .C(n76), .D(regg[115]), .Y(n194) );
  AOI22X1 U317 ( .A(n84), .B(regg[99]), .C(regg[83]), .D(n59), .Y(n195) );
  AOI22X1 U319 ( .A(n84), .B(regg[83]), .C(regg[67]), .D(n51), .Y(n196) );
  AOI22X1 U321 ( .A(n84), .B(regg[67]), .C(regg[51]), .D(n58), .Y(n197) );
  AOI22X1 U323 ( .A(n84), .B(regg[51]), .C(regg[35]), .D(n58), .Y(n198) );
  OAI22X1 U324 ( .A(n64), .B(n795), .C(n794), .D(n73), .Y(n468) );
  OAI22X1 U326 ( .A(n793), .B(n79), .C(n62), .D(n794), .Y(n469) );
  OAI21X1 U328 ( .A(n65), .B(n793), .C(n202), .Y(n470) );
  NAND2X1 U329 ( .A(databus_out[3]), .B(n65), .Y(n202) );
  AOI22X1 U332 ( .A(n85), .B(regg[244]), .C(regg[228]), .D(n51), .Y(n203) );
  AOI22X1 U334 ( .A(n85), .B(regg[228]), .C(regg[212]), .D(n51), .Y(n204) );
  AOI22X1 U336 ( .A(n86), .B(regg[212]), .C(regg[196]), .D(n51), .Y(n205) );
  AOI22X1 U338 ( .A(n86), .B(regg[196]), .C(regg[180]), .D(n52), .Y(n206) );
  AOI22X1 U340 ( .A(n86), .B(regg[180]), .C(regg[164]), .D(n57), .Y(n207) );
  AOI22X1 U342 ( .A(n86), .B(regg[164]), .C(regg[148]), .D(n52), .Y(n208) );
  AOI22X1 U344 ( .A(n87), .B(regg[148]), .C(regg[132]), .D(n52), .Y(n209) );
  AOI22X1 U346 ( .A(n87), .B(regg[132]), .C(regg[116]), .D(n52), .Y(n210) );
  AOI22X1 U348 ( .A(n87), .B(regg[116]), .C(regg[100]), .D(n52), .Y(n211) );
  AOI22X1 U350 ( .A(regg[84]), .B(n61), .C(n76), .D(regg[100]), .Y(n212) );
  AOI22X1 U352 ( .A(n87), .B(regg[84]), .C(regg[68]), .D(n52), .Y(n213) );
  AOI22X1 U354 ( .A(n88), .B(regg[68]), .C(regg[52]), .D(n56), .Y(n214) );
  AOI22X1 U356 ( .A(n88), .B(regg[52]), .C(regg[36]), .D(n56), .Y(n215) );
  OAI22X1 U357 ( .A(n63), .B(n792), .C(n791), .D(n73), .Y(n484) );
  OAI22X1 U359 ( .A(n790), .B(n79), .C(n62), .D(n791), .Y(n485) );
  OAI21X1 U361 ( .A(n65), .B(n790), .C(n219), .Y(n486) );
  NAND2X1 U362 ( .A(databus_out[4]), .B(n63), .Y(n219) );
  AOI22X1 U365 ( .A(n89), .B(regg[245]), .C(regg[229]), .D(n52), .Y(n220) );
  AOI22X1 U367 ( .A(n89), .B(regg[229]), .C(regg[213]), .D(n56), .Y(n221) );
  AOI22X1 U369 ( .A(n89), .B(regg[213]), .C(regg[197]), .D(n53), .Y(n222) );
  AOI22X1 U371 ( .A(n90), .B(regg[197]), .C(regg[181]), .D(n53), .Y(n223) );
  AOI22X1 U373 ( .A(n90), .B(regg[181]), .C(regg[165]), .D(n53), .Y(n224) );
  AOI22X1 U375 ( .A(n90), .B(regg[165]), .C(regg[149]), .D(n53), .Y(n225) );
  AOI22X1 U377 ( .A(n90), .B(regg[149]), .C(regg[133]), .D(n53), .Y(n226) );
  AOI22X1 U379 ( .A(n90), .B(regg[133]), .C(regg[117]), .D(n53), .Y(n227) );
  AOI22X1 U381 ( .A(n91), .B(regg[117]), .C(regg[101]), .D(n55), .Y(n228) );
  AOI22X1 U383 ( .A(regg[85]), .B(n61), .C(n75), .D(regg[101]), .Y(n229) );
  AOI22X1 U385 ( .A(n91), .B(regg[85]), .C(regg[69]), .D(n55), .Y(n230) );
  AOI22X1 U387 ( .A(n92), .B(regg[69]), .C(regg[53]), .D(n55), .Y(n231) );
  AOI22X1 U389 ( .A(n92), .B(regg[53]), .C(regg[37]), .D(n55), .Y(n232) );
  OAI22X1 U390 ( .A(n63), .B(n789), .C(n788), .D(n70), .Y(n500) );
  OAI22X1 U392 ( .A(n787), .B(n78), .C(n62), .D(n788), .Y(n501) );
  OAI21X1 U394 ( .A(n64), .B(n787), .C(n236), .Y(n502) );
  NAND2X1 U395 ( .A(databus_out[5]), .B(n65), .Y(n236) );
  AOI22X1 U398 ( .A(n93), .B(regg[246]), .C(regg[230]), .D(n54), .Y(n237) );
  AOI22X1 U400 ( .A(n93), .B(regg[230]), .C(regg[214]), .D(n54), .Y(n238) );
  AOI22X1 U402 ( .A(n93), .B(regg[214]), .C(regg[198]), .D(n54), .Y(n239) );
  AOI22X1 U404 ( .A(n93), .B(regg[198]), .C(regg[182]), .D(n54), .Y(n240) );
  AOI22X1 U406 ( .A(n93), .B(regg[182]), .C(regg[166]), .D(n54), .Y(n241) );
  AOI22X1 U408 ( .A(n94), .B(regg[166]), .C(regg[150]), .D(n54), .Y(n242) );
  AOI22X1 U410 ( .A(n94), .B(regg[150]), .C(regg[134]), .D(n54), .Y(n243) );
  AOI22X1 U412 ( .A(n94), .B(regg[134]), .C(regg[118]), .D(n53), .Y(n244) );
  AOI22X1 U414 ( .A(n95), .B(regg[118]), .C(regg[102]), .D(n53), .Y(n245) );
  AOI22X1 U416 ( .A(regg[86]), .B(n61), .C(n74), .D(regg[102]), .Y(n246) );
  AOI22X1 U418 ( .A(n95), .B(regg[86]), .C(regg[70]), .D(n53), .Y(n247) );
  AOI22X1 U420 ( .A(n95), .B(regg[70]), .C(regg[54]), .D(n52), .Y(n248) );
  AOI22X1 U422 ( .A(n96), .B(regg[54]), .C(regg[38]), .D(n52), .Y(n249) );
  OAI22X1 U423 ( .A(n63), .B(n786), .C(n785), .D(n70), .Y(n516) );
  OAI22X1 U425 ( .A(n784), .B(n78), .C(n62), .D(n785), .Y(n517) );
  OAI21X1 U427 ( .A(n64), .B(n784), .C(n253), .Y(n518) );
  NAND2X1 U428 ( .A(databus_out[6]), .B(n64), .Y(n253) );
  AOI22X1 U431 ( .A(n89), .B(regg[247]), .C(regg[231]), .D(n51), .Y(n254) );
  AOI22X1 U433 ( .A(n133), .B(regg[231]), .C(regg[215]), .D(n51), .Y(n255) );
  AOI22X1 U435 ( .A(n117), .B(regg[215]), .C(regg[199]), .D(n51), .Y(n256) );
  AOI22X1 U437 ( .A(n117), .B(regg[199]), .C(regg[183]), .D(n51), .Y(n257) );
  AOI22X1 U439 ( .A(n117), .B(regg[183]), .C(regg[167]), .D(n50), .Y(n258) );
  AOI22X1 U441 ( .A(n117), .B(regg[167]), .C(regg[151]), .D(n50), .Y(n259) );
  AOI22X1 U443 ( .A(n117), .B(regg[151]), .C(regg[135]), .D(n50), .Y(n260) );
  AOI22X1 U445 ( .A(n116), .B(regg[135]), .C(regg[119]), .D(n50), .Y(n261) );
  AOI22X1 U447 ( .A(n116), .B(regg[119]), .C(regg[103]), .D(n50), .Y(n262) );
  AOI22X1 U449 ( .A(regg[87]), .B(n61), .C(n76), .D(regg[103]), .Y(n263) );
  AOI22X1 U451 ( .A(n116), .B(regg[87]), .C(regg[71]), .D(n49), .Y(n264) );
  AOI22X1 U453 ( .A(n116), .B(regg[71]), .C(regg[55]), .D(n49), .Y(n265) );
  AOI22X1 U455 ( .A(n116), .B(regg[55]), .C(regg[39]), .D(n49), .Y(n266) );
  OAI22X1 U456 ( .A(n62), .B(n783), .C(n782), .D(n71), .Y(n532) );
  OAI22X1 U458 ( .A(n781), .B(n78), .C(n62), .D(n782), .Y(n533) );
  OAI21X1 U460 ( .A(n65), .B(n781), .C(n270), .Y(n534) );
  NAND2X1 U461 ( .A(databus_out[7]), .B(n65), .Y(n270) );
  AOI22X1 U464 ( .A(n115), .B(regg[248]), .C(regg[232]), .D(n48), .Y(n271) );
  AOI22X1 U466 ( .A(n115), .B(regg[232]), .C(regg[216]), .D(n48), .Y(n272) );
  AOI22X1 U468 ( .A(n115), .B(regg[216]), .C(regg[200]), .D(n48), .Y(n273) );
  AOI22X1 U470 ( .A(n115), .B(regg[200]), .C(regg[184]), .D(n47), .Y(n274) );
  AOI22X1 U472 ( .A(n115), .B(regg[184]), .C(regg[168]), .D(n47), .Y(n275) );
  AOI22X1 U474 ( .A(n114), .B(regg[168]), .C(regg[152]), .D(n47), .Y(n276) );
  AOI22X1 U476 ( .A(n114), .B(regg[152]), .C(regg[136]), .D(n46), .Y(n277) );
  AOI22X1 U478 ( .A(n114), .B(regg[136]), .C(regg[120]), .D(n46), .Y(n278) );
  AOI22X1 U480 ( .A(n114), .B(regg[120]), .C(regg[104]), .D(n46), .Y(n279) );
  AOI22X1 U482 ( .A(regg[88]), .B(n60), .C(n75), .D(regg[104]), .Y(n280) );
  AOI22X1 U484 ( .A(n114), .B(regg[88]), .C(regg[72]), .D(n57), .Y(n281) );
  AOI22X1 U486 ( .A(n113), .B(regg[72]), .C(regg[56]), .D(n57), .Y(n282) );
  AOI22X1 U488 ( .A(n113), .B(regg[56]), .C(regg[40]), .D(n57), .Y(n283) );
  OAI22X1 U489 ( .A(n64), .B(n780), .C(n779), .D(n72), .Y(n548) );
  OAI22X1 U491 ( .A(n778), .B(n79), .C(n62), .D(n779), .Y(n549) );
  OAI21X1 U493 ( .A(n65), .B(n778), .C(n287), .Y(n550) );
  NAND2X1 U494 ( .A(databus_out[8]), .B(n65), .Y(n287) );
  AOI22X1 U497 ( .A(n113), .B(regg[249]), .C(regg[233]), .D(n58), .Y(n288) );
  AOI22X1 U499 ( .A(n113), .B(regg[233]), .C(regg[217]), .D(n60), .Y(n289) );
  AOI22X1 U501 ( .A(n113), .B(regg[217]), .C(regg[201]), .D(n58), .Y(n290) );
  AOI22X1 U503 ( .A(n112), .B(regg[201]), .C(regg[185]), .D(n58), .Y(n291) );
  AOI22X1 U505 ( .A(n112), .B(regg[185]), .C(regg[169]), .D(n58), .Y(n292) );
  AOI22X1 U507 ( .A(n112), .B(regg[169]), .C(regg[153]), .D(n58), .Y(n293) );
  AOI22X1 U509 ( .A(n112), .B(regg[153]), .C(regg[137]), .D(n59), .Y(n294) );
  AOI22X1 U511 ( .A(n112), .B(regg[137]), .C(regg[121]), .D(n59), .Y(n295) );
  AOI22X1 U513 ( .A(n111), .B(regg[121]), .C(regg[105]), .D(n58), .Y(n296) );
  AOI22X1 U515 ( .A(regg[89]), .B(n61), .C(n76), .D(regg[105]), .Y(n297) );
  AOI22X1 U517 ( .A(n111), .B(regg[89]), .C(regg[73]), .D(n59), .Y(n298) );
  AOI22X1 U519 ( .A(n111), .B(regg[73]), .C(regg[57]), .D(n59), .Y(n299) );
  AOI22X1 U521 ( .A(n111), .B(regg[57]), .C(regg[41]), .D(n59), .Y(n300) );
  OAI22X1 U522 ( .A(n64), .B(n777), .C(n776), .D(n72), .Y(n564) );
  OAI22X1 U524 ( .A(n775), .B(n78), .C(n62), .D(n776), .Y(n565) );
  OAI21X1 U526 ( .A(n65), .B(n775), .C(n304), .Y(n566) );
  NAND2X1 U527 ( .A(databus_out[9]), .B(n62), .Y(n304) );
  AOI22X1 U530 ( .A(n111), .B(regg[250]), .C(regg[234]), .D(n57), .Y(n305) );
  AOI22X1 U532 ( .A(n110), .B(regg[234]), .C(regg[218]), .D(n57), .Y(n306) );
  AOI22X1 U534 ( .A(n110), .B(regg[218]), .C(regg[202]), .D(n57), .Y(n307) );
  AOI22X1 U536 ( .A(n110), .B(regg[202]), .C(regg[186]), .D(n56), .Y(n308) );
  AOI22X1 U538 ( .A(n110), .B(regg[186]), .C(regg[170]), .D(n56), .Y(n309) );
  AOI22X1 U540 ( .A(n110), .B(regg[170]), .C(regg[154]), .D(n56), .Y(n310) );
  AOI22X1 U542 ( .A(n109), .B(regg[154]), .C(regg[138]), .D(n56), .Y(n311) );
  AOI22X1 U544 ( .A(n109), .B(regg[138]), .C(regg[122]), .D(n56), .Y(n312) );
  AOI22X1 U546 ( .A(n109), .B(regg[122]), .C(regg[106]), .D(n56), .Y(n313) );
  AOI22X1 U548 ( .A(regg[90]), .B(n61), .C(n75), .D(regg[106]), .Y(n314) );
  AOI22X1 U550 ( .A(n109), .B(regg[90]), .C(regg[74]), .D(n55), .Y(n315) );
  AOI22X1 U552 ( .A(n109), .B(regg[74]), .C(regg[58]), .D(n55), .Y(n316) );
  AOI22X1 U554 ( .A(n108), .B(regg[58]), .C(regg[42]), .D(n55), .Y(n317) );
  OAI22X1 U555 ( .A(n63), .B(n774), .C(n773), .D(n72), .Y(n580) );
  OAI22X1 U557 ( .A(n63), .B(n773), .C(n772), .D(n74), .Y(n581) );
  OAI21X1 U559 ( .A(n64), .B(n772), .C(n321), .Y(n582) );
  NAND2X1 U560 ( .A(databus_out[10]), .B(n61), .Y(n321) );
  AOI22X1 U563 ( .A(n108), .B(regg[251]), .C(regg[235]), .D(n54), .Y(n322) );
  AOI22X1 U565 ( .A(n108), .B(regg[235]), .C(regg[219]), .D(n54), .Y(n323) );
  AOI22X1 U567 ( .A(n108), .B(regg[219]), .C(regg[203]), .D(n54), .Y(n324) );
  AOI22X1 U569 ( .A(n108), .B(regg[203]), .C(regg[187]), .D(n54), .Y(n325) );
  AOI22X1 U571 ( .A(n107), .B(regg[187]), .C(regg[171]), .D(n53), .Y(n326) );
  AOI22X1 U573 ( .A(n107), .B(regg[171]), .C(regg[155]), .D(n53), .Y(n327) );
  AOI22X1 U575 ( .A(n107), .B(regg[155]), .C(regg[139]), .D(n52), .Y(n328) );
  AOI22X1 U577 ( .A(n107), .B(regg[139]), .C(regg[123]), .D(n52), .Y(n329) );
  AOI22X1 U579 ( .A(n106), .B(regg[123]), .C(regg[107]), .D(n51), .Y(n330) );
  AOI22X1 U581 ( .A(regg[91]), .B(n61), .C(n77), .D(regg[107]), .Y(n331) );
  AOI22X1 U583 ( .A(n106), .B(regg[91]), .C(regg[75]), .D(n51), .Y(n332) );
  AOI22X1 U585 ( .A(n106), .B(regg[75]), .C(regg[59]), .D(n50), .Y(n333) );
  AOI22X1 U587 ( .A(n106), .B(regg[59]), .C(regg[43]), .D(n50), .Y(n334) );
  OAI22X1 U588 ( .A(n63), .B(n771), .C(n770), .D(n74), .Y(n596) );
  OAI22X1 U590 ( .A(n63), .B(n770), .C(n769), .D(n73), .Y(n597) );
  OAI21X1 U592 ( .A(n64), .B(n769), .C(n338), .Y(n598) );
  NAND2X1 U593 ( .A(databus_out[11]), .B(n63), .Y(n338) );
  AOI22X1 U596 ( .A(n106), .B(regg[252]), .C(regg[236]), .D(n48), .Y(n339) );
  AOI22X1 U598 ( .A(n105), .B(regg[236]), .C(regg[220]), .D(n47), .Y(n340) );
  AOI22X1 U600 ( .A(n105), .B(regg[220]), .C(regg[204]), .D(n47), .Y(n341) );
  AOI22X1 U602 ( .A(n105), .B(regg[204]), .C(regg[188]), .D(n46), .Y(n342) );
  AOI22X1 U604 ( .A(n105), .B(regg[188]), .C(regg[172]), .D(n46), .Y(n343) );
  AOI22X1 U606 ( .A(n105), .B(regg[172]), .C(regg[156]), .D(n60), .Y(n344) );
  AOI22X1 U608 ( .A(n104), .B(regg[156]), .C(regg[140]), .D(n60), .Y(n345) );
  AOI22X1 U610 ( .A(n104), .B(regg[140]), .C(regg[124]), .D(n60), .Y(n346) );
  AOI22X1 U612 ( .A(n104), .B(regg[124]), .C(regg[108]), .D(n60), .Y(n347) );
  AOI22X1 U614 ( .A(regg[92]), .B(n61), .C(n77), .D(regg[108]), .Y(n348) );
  AOI22X1 U616 ( .A(n104), .B(regg[92]), .C(regg[76]), .D(n60), .Y(n349) );
  AOI22X1 U618 ( .A(n104), .B(regg[76]), .C(regg[60]), .D(n59), .Y(n350) );
  AOI22X1 U620 ( .A(n103), .B(regg[60]), .C(regg[44]), .D(n59), .Y(n351) );
  OAI22X1 U621 ( .A(n63), .B(n768), .C(n767), .D(n74), .Y(n612) );
  OAI22X1 U623 ( .A(n63), .B(n767), .C(n766), .D(n71), .Y(n613) );
  OAI21X1 U625 ( .A(n64), .B(n766), .C(n355), .Y(n614) );
  NAND2X1 U626 ( .A(databus_out[12]), .B(n62), .Y(n355) );
  AOI22X1 U629 ( .A(n103), .B(regg[253]), .C(regg[237]), .D(n57), .Y(n356) );
  AOI22X1 U631 ( .A(n103), .B(regg[237]), .C(regg[221]), .D(n57), .Y(n357) );
  AOI22X1 U633 ( .A(n103), .B(regg[221]), .C(regg[205]), .D(n56), .Y(n358) );
  AOI22X1 U635 ( .A(n103), .B(regg[205]), .C(regg[189]), .D(n56), .Y(n359) );
  AOI22X1 U637 ( .A(n102), .B(regg[189]), .C(regg[173]), .D(n56), .Y(n360) );
  AOI22X1 U639 ( .A(n102), .B(regg[173]), .C(regg[157]), .D(n55), .Y(n361) );
  AOI22X1 U641 ( .A(n102), .B(regg[157]), .C(regg[141]), .D(n55), .Y(n362) );
  AOI22X1 U643 ( .A(n102), .B(regg[141]), .C(regg[125]), .D(n55), .Y(n363) );
  AOI22X1 U645 ( .A(n102), .B(regg[125]), .C(regg[109]), .D(n54), .Y(n364) );
  AOI22X1 U647 ( .A(regg[93]), .B(n61), .C(n77), .D(regg[109]), .Y(n365) );
  AOI22X1 U649 ( .A(n101), .B(regg[93]), .C(regg[77]), .D(n53), .Y(n366) );
  AOI22X1 U651 ( .A(n101), .B(regg[77]), .C(regg[61]), .D(n53), .Y(n367) );
  AOI22X1 U653 ( .A(n101), .B(regg[61]), .C(regg[45]), .D(n52), .Y(n368) );
  OAI22X1 U654 ( .A(n64), .B(n765), .C(n764), .D(n72), .Y(n628) );
  OAI22X1 U656 ( .A(n63), .B(n764), .C(n763), .D(n71), .Y(n629) );
  OAI21X1 U658 ( .A(n65), .B(n763), .C(n372), .Y(n630) );
  NAND2X1 U659 ( .A(databus_out[13]), .B(n65), .Y(n372) );
  AOI22X1 U662 ( .A(n101), .B(regg[254]), .C(regg[238]), .D(n48), .Y(n373) );
  AOI22X1 U664 ( .A(n101), .B(regg[238]), .C(regg[222]), .D(n47), .Y(n374) );
  AOI22X1 U666 ( .A(n100), .B(regg[222]), .C(regg[206]), .D(n46), .Y(n375) );
  AOI22X1 U668 ( .A(n100), .B(regg[206]), .C(regg[190]), .D(n60), .Y(n376) );
  AOI22X1 U670 ( .A(n100), .B(regg[190]), .C(regg[174]), .D(n60), .Y(n377) );
  AOI22X1 U672 ( .A(n100), .B(regg[174]), .C(regg[158]), .D(n60), .Y(n378) );
  AOI22X1 U674 ( .A(n100), .B(regg[158]), .C(regg[142]), .D(n59), .Y(n379) );
  AOI22X1 U676 ( .A(n99), .B(regg[142]), .C(regg[126]), .D(n59), .Y(n380) );
  AOI22X1 U678 ( .A(n99), .B(regg[126]), .C(regg[110]), .D(n58), .Y(n381) );
  AOI22X1 U680 ( .A(regg[94]), .B(n61), .C(n76), .D(regg[110]), .Y(n382) );
  AOI22X1 U682 ( .A(n99), .B(regg[94]), .C(regg[78]), .D(n56), .Y(n383) );
  AOI22X1 U684 ( .A(n99), .B(regg[78]), .C(regg[62]), .D(n55), .Y(n384) );
  AOI22X1 U686 ( .A(n99), .B(regg[62]), .C(regg[46]), .D(n55), .Y(n385) );
  OAI22X1 U687 ( .A(n63), .B(n762), .C(n761), .D(n72), .Y(n644) );
  OAI22X1 U689 ( .A(n63), .B(n761), .C(n760), .D(n71), .Y(n645) );
  OAI21X1 U691 ( .A(n65), .B(n760), .C(n389), .Y(n646) );
  NAND2X1 U692 ( .A(databus_out[14]), .B(n65), .Y(n389) );
  AOI22X1 U695 ( .A(n98), .B(regg[255]), .C(regg[239]), .D(n48), .Y(n390) );
  AOI22X1 U697 ( .A(n98), .B(regg[239]), .C(regg[223]), .D(n46), .Y(n391) );
  AOI22X1 U699 ( .A(n98), .B(regg[223]), .C(regg[207]), .D(n50), .Y(n392) );
  AOI22X1 U701 ( .A(n98), .B(regg[207]), .C(regg[191]), .D(n49), .Y(n393) );
  AOI22X1 U703 ( .A(n98), .B(regg[191]), .C(regg[175]), .D(n58), .Y(n394) );
  AOI22X1 U705 ( .A(n97), .B(regg[175]), .C(regg[159]), .D(n49), .Y(n395) );
  AOI22X1 U707 ( .A(n97), .B(regg[159]), .C(regg[143]), .D(n55), .Y(n396) );
  AOI22X1 U709 ( .A(n97), .B(regg[143]), .C(regg[127]), .D(n57), .Y(n397) );
  AOI22X1 U711 ( .A(n97), .B(regg[127]), .C(regg[111]), .D(n60), .Y(n398) );
  AOI22X1 U713 ( .A(regg[95]), .B(n61), .C(n75), .D(regg[111]), .Y(n399) );
  AOI22X1 U715 ( .A(n97), .B(regg[95]), .C(regg[79]), .D(n51), .Y(n400) );
  AOI22X1 U717 ( .A(n107), .B(regg[79]), .C(regg[63]), .D(n54), .Y(n401) );
  AOI22X1 U719 ( .A(n96), .B(regg[63]), .C(regg[47]), .D(n52), .Y(n402) );
  OAI22X1 U720 ( .A(n64), .B(n759), .C(n758), .D(n70), .Y(n660) );
  OAI22X1 U722 ( .A(n62), .B(n758), .C(n757), .D(n70), .Y(n661) );
  OAI21X1 U725 ( .A(n65), .B(n757), .C(n406), .Y(n662) );
  NAND2X1 U726 ( .A(databus_out[15]), .B(n65), .Y(n406) );
  INVX1 U2 ( .A(n150), .Y(n1) );
  BUFX2 U3 ( .A(n37), .Y(n2) );
  BUFX2 U4 ( .A(n17), .Y(n37) );
  BUFX4 U5 ( .A(n14), .Y(n4) );
  BUFX2 U6 ( .A(n12), .Y(n3) );
  BUFX2 U7 ( .A(n10), .Y(n38) );
  BUFX4 U8 ( .A(n519), .Y(n44) );
  BUFX4 U9 ( .A(n10), .Y(n39) );
  BUFX2 U10 ( .A(n14), .Y(n16) );
  INVX2 U11 ( .A(n15), .Y(n17) );
  BUFX4 U12 ( .A(n12), .Y(n9) );
  INVX2 U13 ( .A(n167), .Y(n515) );
  INVX4 U14 ( .A(n16), .Y(n11) );
  BUFX4 U15 ( .A(n514), .Y(n36) );
  INVX2 U16 ( .A(n6), .Y(n5) );
  INVX4 U17 ( .A(n36), .Y(n6) );
  BUFX2 U18 ( .A(n44), .Y(n41) );
  BUFX2 U19 ( .A(n35), .Y(n34) );
  INVX8 U20 ( .A(n6), .Y(n7) );
  INVX8 U21 ( .A(n6), .Y(n8) );
  INVX2 U22 ( .A(n167), .Y(n10) );
  BUFX4 U23 ( .A(n515), .Y(n19) );
  INVX8 U24 ( .A(n11), .Y(n12) );
  INVX1 U25 ( .A(n150), .Y(n13) );
  INVX4 U26 ( .A(n150), .Y(n514) );
  BUFX2 U27 ( .A(n42), .Y(n45) );
  INVX2 U28 ( .A(n15), .Y(n14) );
  INVX2 U29 ( .A(n166), .Y(n32) );
  NAND2X1 U30 ( .A(row_sel[0]), .B(row_sel[1]), .Y(n15) );
  INVX2 U31 ( .A(n68), .Y(n53) );
  INVX2 U32 ( .A(n69), .Y(n47) );
  INVX2 U33 ( .A(n68), .Y(n56) );
  INVX2 U34 ( .A(n69), .Y(n48) );
  INVX2 U35 ( .A(n69), .Y(n50) );
  INVX2 U36 ( .A(n69), .Y(n49) );
  INVX2 U37 ( .A(n68), .Y(n55) );
  INVX2 U38 ( .A(n69), .Y(n51) );
  INVX2 U39 ( .A(n68), .Y(n54) );
  INVX2 U40 ( .A(n68), .Y(n52) );
  INVX2 U41 ( .A(n67), .Y(n59) );
  INVX2 U42 ( .A(n67), .Y(n58) );
  INVX2 U43 ( .A(n67), .Y(n57) );
  INVX2 U44 ( .A(n67), .Y(n60) );
  INVX2 U45 ( .A(n67), .Y(n61) );
  INVX2 U46 ( .A(n66), .Y(n62) );
  INVX2 U47 ( .A(n66), .Y(n63) );
  INVX2 U48 ( .A(n66), .Y(n64) );
  INVX2 U49 ( .A(n66), .Y(n65) );
  INVX2 U50 ( .A(n70), .Y(n46) );
  BUFX2 U51 ( .A(n135), .Y(n69) );
  BUFX2 U52 ( .A(n135), .Y(n68) );
  BUFX2 U53 ( .A(n148), .Y(n67) );
  BUFX2 U54 ( .A(n148), .Y(n66) );
  BUFX2 U55 ( .A(n135), .Y(n70) );
  BUFX2 U56 ( .A(n133), .Y(n73) );
  BUFX2 U57 ( .A(n133), .Y(n72) );
  BUFX2 U58 ( .A(n133), .Y(n71) );
  BUFX2 U59 ( .A(n132), .Y(n74) );
  BUFX2 U60 ( .A(n131), .Y(n77) );
  BUFX2 U61 ( .A(n132), .Y(n76) );
  BUFX2 U62 ( .A(n132), .Y(n75) );
  BUFX2 U63 ( .A(n131), .Y(n78) );
  BUFX2 U64 ( .A(n131), .Y(n79) );
  BUFX2 U65 ( .A(n130), .Y(n80) );
  BUFX2 U66 ( .A(n130), .Y(n81) );
  BUFX2 U67 ( .A(n130), .Y(n82) );
  BUFX2 U68 ( .A(n129), .Y(n83) );
  BUFX2 U69 ( .A(n129), .Y(n84) );
  BUFX2 U70 ( .A(n129), .Y(n85) );
  BUFX2 U71 ( .A(n128), .Y(n86) );
  BUFX2 U72 ( .A(n128), .Y(n87) );
  BUFX2 U73 ( .A(n128), .Y(n88) );
  BUFX2 U74 ( .A(n127), .Y(n90) );
  BUFX2 U75 ( .A(n127), .Y(n91) );
  BUFX2 U76 ( .A(n126), .Y(n92) );
  BUFX2 U77 ( .A(n126), .Y(n93) );
  BUFX2 U78 ( .A(n126), .Y(n94) );
  BUFX2 U79 ( .A(n125), .Y(n95) );
  BUFX2 U80 ( .A(n127), .Y(n89) );
  BUFX2 U81 ( .A(n118), .Y(n117) );
  BUFX2 U82 ( .A(n118), .Y(n116) );
  BUFX2 U83 ( .A(n119), .Y(n115) );
  BUFX2 U84 ( .A(n119), .Y(n114) );
  BUFX2 U85 ( .A(n119), .Y(n113) );
  BUFX2 U86 ( .A(n120), .Y(n112) );
  BUFX2 U87 ( .A(n120), .Y(n111) );
  BUFX2 U88 ( .A(n120), .Y(n110) );
  BUFX2 U89 ( .A(n121), .Y(n109) );
  BUFX2 U90 ( .A(n121), .Y(n108) );
  BUFX2 U91 ( .A(n122), .Y(n106) );
  BUFX2 U92 ( .A(n122), .Y(n105) );
  BUFX2 U93 ( .A(n122), .Y(n104) );
  BUFX2 U94 ( .A(n123), .Y(n103) );
  BUFX2 U95 ( .A(n123), .Y(n102) );
  BUFX2 U96 ( .A(n123), .Y(n101) );
  BUFX2 U97 ( .A(n124), .Y(n100) );
  BUFX2 U98 ( .A(n124), .Y(n99) );
  BUFX2 U99 ( .A(n124), .Y(n98) );
  BUFX2 U100 ( .A(n125), .Y(n97) );
  BUFX2 U101 ( .A(n121), .Y(n107) );
  BUFX2 U102 ( .A(n125), .Y(n96) );
  BUFX2 U103 ( .A(n149), .Y(n135) );
  BUFX2 U104 ( .A(n149), .Y(n148) );
  BUFX2 U105 ( .A(n149), .Y(n118) );
  BUFX2 U106 ( .A(n149), .Y(n119) );
  BUFX2 U107 ( .A(n118), .Y(n120) );
  BUFX2 U108 ( .A(n149), .Y(n130) );
  BUFX2 U109 ( .A(n149), .Y(n129) );
  BUFX2 U110 ( .A(n149), .Y(n128) );
  BUFX2 U111 ( .A(n149), .Y(n126) );
  BUFX2 U112 ( .A(n149), .Y(n127) );
  BUFX2 U113 ( .A(n119), .Y(n122) );
  BUFX2 U114 ( .A(n123), .Y(n131) );
  BUFX2 U115 ( .A(n130), .Y(n123) );
  BUFX2 U116 ( .A(n129), .Y(n124) );
  BUFX2 U117 ( .A(n122), .Y(n132) );
  BUFX2 U118 ( .A(n128), .Y(n121) );
  BUFX2 U119 ( .A(n126), .Y(n125) );
  BUFX2 U120 ( .A(n120), .Y(n133) );
  INVX2 U121 ( .A(strb_matrix), .Y(n149) );
  BUFX2 U122 ( .A(n514), .Y(n35) );
  BUFX2 U123 ( .A(n39), .Y(n18) );
  BUFX2 U124 ( .A(n38), .Y(n20) );
  BUFX2 U125 ( .A(n38), .Y(n21) );
  BUFX2 U126 ( .A(n40), .Y(n22) );
  BUFX2 U127 ( .A(n40), .Y(n23) );
  BUFX2 U128 ( .A(n40), .Y(n24) );
  BUFX2 U129 ( .A(n39), .Y(n25) );
  BUFX2 U130 ( .A(n39), .Y(n26) );
  BUFX2 U131 ( .A(n38), .Y(n27) );
  BUFX2 U132 ( .A(n38), .Y(n28) );
  BUFX2 U133 ( .A(n38), .Y(n29) );
  BUFX2 U134 ( .A(n38), .Y(n30) );
  BUFX2 U135 ( .A(n38), .Y(n31) );
  BUFX2 U136 ( .A(n38), .Y(n40) );
  INVX2 U137 ( .A(n166), .Y(n519) );
  BUFX2 U138 ( .A(n32), .Y(n42) );
  BUFX4 U139 ( .A(n13), .Y(n33) );
  BUFX4 U140 ( .A(n519), .Y(n43) );
  INVX2 U141 ( .A(row_sel[1]), .Y(n165) );
  OR2X2 U142 ( .A(row_sel[0]), .B(n165), .Y(n150) );
  AOI22X1 U143 ( .A(regg[0]), .B(n9), .C(regg[64]), .D(n33), .Y(n183) );
  NAND2X1 U144 ( .A(n165), .B(row_sel[0]), .Y(n166) );
  OR2X2 U145 ( .A(row_sel[0]), .B(row_sel[1]), .Y(n167) );
  AOI22X1 U146 ( .A(regg[128]), .B(n43), .C(regg[192]), .D(n20), .Y(n182) );
  NAND2X1 U147 ( .A(n183), .B(n182), .Y(row[0]) );
  AOI22X1 U148 ( .A(regg[1]), .B(n2), .C(regg[65]), .D(n8), .Y(n199) );
  AOI22X1 U149 ( .A(regg[129]), .B(n43), .C(regg[193]), .D(n19), .Y(n184) );
  NAND2X1 U150 ( .A(n199), .B(n184), .Y(row[1]) );
  AOI22X1 U151 ( .A(regg[2]), .B(n3), .C(regg[66]), .D(n34), .Y(n201) );
  AOI22X1 U152 ( .A(regg[130]), .B(n41), .C(regg[194]), .D(n30), .Y(n200) );
  NAND2X1 U153 ( .A(n201), .B(n200), .Y(row[2]) );
  AOI22X1 U154 ( .A(regg[3]), .B(n9), .C(regg[67]), .D(n7), .Y(n217) );
  AOI22X1 U155 ( .A(regg[131]), .B(n45), .C(regg[195]), .D(n21), .Y(n216) );
  NAND2X1 U156 ( .A(n217), .B(n216), .Y(row[3]) );
  AOI22X1 U157 ( .A(regg[4]), .B(n2), .C(regg[68]), .D(n33), .Y(n233) );
  AOI22X1 U158 ( .A(regg[132]), .B(n43), .C(regg[196]), .D(n22), .Y(n218) );
  NAND2X1 U159 ( .A(n233), .B(n218), .Y(row[4]) );
  AOI22X1 U160 ( .A(regg[5]), .B(n3), .C(regg[69]), .D(n8), .Y(n235) );
  AOI22X1 U161 ( .A(regg[133]), .B(n43), .C(regg[197]), .D(n30), .Y(n234) );
  NAND2X1 U162 ( .A(n235), .B(n234), .Y(row[5]) );
  AOI22X1 U163 ( .A(regg[6]), .B(n9), .C(regg[70]), .D(n33), .Y(n251) );
  AOI22X1 U164 ( .A(regg[134]), .B(n41), .C(regg[198]), .D(n23), .Y(n250) );
  NAND2X1 U165 ( .A(n251), .B(n250), .Y(row[6]) );
  AOI22X1 U166 ( .A(regg[7]), .B(n9), .C(regg[71]), .D(n7), .Y(n267) );
  AOI22X1 U167 ( .A(regg[135]), .B(n45), .C(regg[199]), .D(n24), .Y(n252) );
  NAND2X1 U168 ( .A(n267), .B(n252), .Y(row[7]) );
  AOI22X1 U169 ( .A(regg[8]), .B(n2), .C(regg[72]), .D(n34), .Y(n269) );
  AOI22X1 U170 ( .A(regg[136]), .B(n43), .C(regg[200]), .D(n30), .Y(n268) );
  NAND2X1 U171 ( .A(n269), .B(n268), .Y(row[8]) );
  AOI22X1 U172 ( .A(regg[9]), .B(n9), .C(regg[73]), .D(n33), .Y(n285) );
  AOI22X1 U173 ( .A(regg[137]), .B(n41), .C(regg[201]), .D(n30), .Y(n284) );
  NAND2X1 U174 ( .A(n285), .B(n284), .Y(row[9]) );
  AOI22X1 U175 ( .A(regg[10]), .B(n3), .C(regg[74]), .D(n8), .Y(n301) );
  AOI22X1 U176 ( .A(regg[138]), .B(n43), .C(regg[202]), .D(n30), .Y(n286) );
  NAND2X1 U177 ( .A(n301), .B(n286), .Y(row[10]) );
  AOI22X1 U178 ( .A(regg[11]), .B(n9), .C(regg[75]), .D(n7), .Y(n303) );
  AOI22X1 U179 ( .A(regg[139]), .B(n43), .C(regg[203]), .D(n25), .Y(n302) );
  NAND2X1 U180 ( .A(n303), .B(n302), .Y(row[11]) );
  AOI22X1 U181 ( .A(regg[12]), .B(n2), .C(regg[76]), .D(n33), .Y(n319) );
  AOI22X1 U182 ( .A(regg[140]), .B(n45), .C(regg[204]), .D(n26), .Y(n318) );
  NAND2X1 U183 ( .A(n319), .B(n318), .Y(row[12]) );
  AOI22X1 U184 ( .A(regg[13]), .B(n3), .C(regg[77]), .D(n8), .Y(n335) );
  AOI22X1 U185 ( .A(regg[141]), .B(n43), .C(regg[205]), .D(n30), .Y(n320) );
  NAND2X1 U186 ( .A(n335), .B(n320), .Y(row[13]) );
  AOI22X1 U187 ( .A(regg[14]), .B(n3), .C(regg[78]), .D(n34), .Y(n337) );
  AOI22X1 U188 ( .A(regg[142]), .B(n41), .C(regg[206]), .D(n30), .Y(n336) );
  NAND2X1 U189 ( .A(n337), .B(n336), .Y(row[14]) );
  AOI22X1 U190 ( .A(regg[15]), .B(n3), .C(regg[79]), .D(n7), .Y(n353) );
  AOI22X1 U191 ( .A(regg[143]), .B(n45), .C(regg[207]), .D(n30), .Y(n352) );
  NAND2X1 U192 ( .A(n353), .B(n352), .Y(row[15]) );
  NAND2X1 U193 ( .A(n1), .B(regg[80]), .Y(n370) );
  NAND2X1 U194 ( .A(regg[208]), .B(n10), .Y(n369) );
  AOI22X1 U195 ( .A(regg[16]), .B(n17), .C(regg[144]), .D(n519), .Y(n354) );
  NAND3X1 U196 ( .A(n354), .B(n370), .C(n369), .Y(row[16]) );
  AOI22X1 U197 ( .A(n32), .B(regg[145]), .C(regg[17]), .D(n17), .Y(n387) );
  NAND2X1 U198 ( .A(regg[209]), .B(n10), .Y(n386) );
  NAND2X1 U199 ( .A(n1), .B(regg[81]), .Y(n371) );
  NAND3X1 U201 ( .A(n387), .B(n386), .C(n371), .Y(row[17]) );
  AOI22X1 U203 ( .A(regg[18]), .B(n4), .C(regg[82]), .D(n35), .Y(n403) );
  AOI22X1 U205 ( .A(regg[146]), .B(n42), .C(regg[210]), .D(n19), .Y(n388) );
  NAND2X1 U207 ( .A(n403), .B(n388), .Y(row[18]) );
  AOI22X1 U209 ( .A(regg[19]), .B(n37), .C(regg[83]), .D(n33), .Y(n405) );
  AOI22X1 U211 ( .A(regg[147]), .B(n44), .C(regg[211]), .D(n38), .Y(n404) );
  NAND2X1 U213 ( .A(n405), .B(n404), .Y(row[19]) );
  AOI22X1 U215 ( .A(regg[20]), .B(n12), .C(regg[84]), .D(n8), .Y(n408) );
  AOI22X1 U217 ( .A(regg[148]), .B(n43), .C(regg[212]), .D(n21), .Y(n407) );
  NAND2X1 U219 ( .A(n408), .B(n407), .Y(row[20]) );
  AOI22X1 U221 ( .A(regg[21]), .B(n9), .C(regg[85]), .D(n8), .Y(n410) );
  AOI22X1 U223 ( .A(regg[149]), .B(n43), .C(regg[213]), .D(n23), .Y(n409) );
  NAND2X1 U226 ( .A(n410), .B(n409), .Y(row[21]) );
  AOI22X1 U228 ( .A(regg[22]), .B(n12), .C(regg[86]), .D(n7), .Y(n412) );
  AOI22X1 U231 ( .A(regg[150]), .B(n45), .C(regg[214]), .D(n26), .Y(n411) );
  NAND2X1 U232 ( .A(n412), .B(n411), .Y(row[22]) );
  AOI22X1 U234 ( .A(regg[23]), .B(n9), .C(regg[87]), .D(n8), .Y(n414) );
  AOI22X1 U236 ( .A(regg[151]), .B(n41), .C(regg[215]), .D(n25), .Y(n413) );
  NAND2X1 U238 ( .A(n414), .B(n413), .Y(row[23]) );
  AOI22X1 U240 ( .A(regg[24]), .B(n37), .C(regg[88]), .D(n34), .Y(n416) );
  AOI22X1 U242 ( .A(regg[152]), .B(n43), .C(regg[216]), .D(n27), .Y(n415) );
  NAND2X1 U244 ( .A(n416), .B(n415), .Y(row[24]) );
  AOI22X1 U246 ( .A(regg[25]), .B(n9), .C(regg[89]), .D(n8), .Y(n418) );
  AOI22X1 U248 ( .A(regg[153]), .B(n43), .C(regg[217]), .D(n29), .Y(n417) );
  NAND2X1 U250 ( .A(n418), .B(n417), .Y(row[25]) );
  AOI22X1 U252 ( .A(regg[26]), .B(n37), .C(regg[90]), .D(n7), .Y(n423) );
  AOI22X1 U254 ( .A(regg[154]), .B(n43), .C(regg[218]), .D(n31), .Y(n419) );
  NAND2X1 U256 ( .A(n423), .B(n419), .Y(row[26]) );
  AOI22X1 U259 ( .A(regg[27]), .B(n9), .C(regg[91]), .D(n33), .Y(n425) );
  AOI22X1 U261 ( .A(regg[155]), .B(n41), .C(regg[219]), .D(n31), .Y(n424) );
  NAND2X1 U264 ( .A(n425), .B(n424), .Y(row[27]) );
  AOI22X1 U265 ( .A(regg[28]), .B(n3), .C(regg[92]), .D(n7), .Y(n427) );
  AOI22X1 U267 ( .A(regg[156]), .B(n43), .C(regg[220]), .D(n31), .Y(n426) );
  NAND2X1 U269 ( .A(n427), .B(n426), .Y(row[28]) );
  AOI22X1 U271 ( .A(regg[29]), .B(n9), .C(regg[93]), .D(n8), .Y(n429) );
  AOI22X1 U273 ( .A(regg[157]), .B(n43), .C(regg[221]), .D(n30), .Y(n428) );
  NAND2X1 U275 ( .A(n429), .B(n428), .Y(row[29]) );
  AOI22X1 U277 ( .A(regg[30]), .B(n9), .C(regg[94]), .D(n7), .Y(n431) );
  AOI22X1 U279 ( .A(regg[158]), .B(n43), .C(regg[222]), .D(n30), .Y(n430) );
  NAND2X1 U281 ( .A(n431), .B(n430), .Y(row[30]) );
  AOI22X1 U283 ( .A(regg[31]), .B(n3), .C(regg[95]), .D(n8), .Y(n433) );
  AOI22X1 U285 ( .A(regg[159]), .B(n41), .C(regg[223]), .D(n18), .Y(n432) );
  NAND2X1 U287 ( .A(n433), .B(n432), .Y(row[31]) );
  NAND2X1 U289 ( .A(n514), .B(regg[96]), .Y(n439) );
  NAND2X1 U292 ( .A(regg[224]), .B(n10), .Y(n435) );
  AOI22X1 U294 ( .A(regg[32]), .B(n17), .C(regg[160]), .D(n519), .Y(n434) );
  NAND3X1 U297 ( .A(n439), .B(n434), .C(n435), .Y(row[32]) );
  NAND2X1 U298 ( .A(regg[97]), .B(n13), .Y(n442) );
  NAND2X1 U300 ( .A(regg[225]), .B(n10), .Y(n441) );
  AOI22X1 U302 ( .A(regg[33]), .B(n17), .C(regg[161]), .D(n519), .Y(n440) );
  NAND3X1 U304 ( .A(n442), .B(n441), .C(n440), .Y(row[33]) );
  AOI22X1 U306 ( .A(regg[34]), .B(n16), .C(regg[98]), .D(n35), .Y(n444) );
  AOI22X1 U308 ( .A(regg[162]), .B(n42), .C(regg[226]), .D(n39), .Y(n443) );
  NAND2X1 U310 ( .A(n444), .B(n443), .Y(row[34]) );
  AOI22X1 U312 ( .A(regg[35]), .B(n12), .C(regg[99]), .D(n7), .Y(n446) );
  AOI22X1 U314 ( .A(regg[163]), .B(n44), .C(regg[227]), .D(n18), .Y(n445) );
  NAND2X1 U316 ( .A(n446), .B(n445), .Y(row[35]) );
  AOI22X1 U318 ( .A(regg[36]), .B(n12), .C(regg[100]), .D(n34), .Y(n448) );
  AOI22X1 U320 ( .A(regg[164]), .B(n41), .C(regg[228]), .D(n22), .Y(n447) );
  NAND2X1 U322 ( .A(n448), .B(n447), .Y(row[36]) );
  AOI22X1 U325 ( .A(regg[37]), .B(n12), .C(regg[101]), .D(n33), .Y(n450) );
  AOI22X1 U327 ( .A(regg[165]), .B(n43), .C(regg[229]), .D(n24), .Y(n449) );
  NAND2X1 U330 ( .A(n450), .B(n449), .Y(row[37]) );
  AOI22X1 U331 ( .A(regg[38]), .B(n37), .C(regg[102]), .D(n34), .Y(n455) );
  AOI22X1 U333 ( .A(regg[166]), .B(n43), .C(regg[230]), .D(n26), .Y(n451) );
  NAND2X1 U335 ( .A(n455), .B(n451), .Y(row[38]) );
  AOI22X1 U337 ( .A(regg[39]), .B(n12), .C(regg[103]), .D(n7), .Y(n457) );
  AOI22X1 U339 ( .A(regg[167]), .B(n45), .C(regg[231]), .D(n28), .Y(n456) );
  NAND2X1 U341 ( .A(n457), .B(n456), .Y(row[39]) );
  AOI22X1 U343 ( .A(regg[40]), .B(n12), .C(regg[104]), .D(n8), .Y(n459) );
  AOI22X1 U345 ( .A(regg[168]), .B(n41), .C(regg[232]), .D(n27), .Y(n458) );
  NAND2X1 U347 ( .A(n459), .B(n458), .Y(row[40]) );
  AOI22X1 U349 ( .A(regg[41]), .B(n12), .C(regg[105]), .D(n33), .Y(n461) );
  AOI22X1 U351 ( .A(regg[169]), .B(n43), .C(regg[233]), .D(n29), .Y(n460) );
  NAND2X1 U353 ( .A(n461), .B(n460), .Y(row[41]) );
  AOI22X1 U355 ( .A(regg[42]), .B(n12), .C(regg[106]), .D(n34), .Y(n463) );
  AOI22X1 U358 ( .A(regg[170]), .B(n45), .C(regg[234]), .D(n27), .Y(n462) );
  NAND2X1 U360 ( .A(n463), .B(n462), .Y(row[42]) );
  AOI22X1 U363 ( .A(regg[43]), .B(n3), .C(regg[107]), .D(n8), .Y(n465) );
  AOI22X1 U364 ( .A(regg[171]), .B(n43), .C(regg[235]), .D(n29), .Y(n464) );
  NAND2X1 U366 ( .A(n465), .B(n464), .Y(row[43]) );
  AOI22X1 U368 ( .A(regg[44]), .B(n2), .C(regg[108]), .D(n33), .Y(n467) );
  AOI22X1 U370 ( .A(regg[172]), .B(n43), .C(regg[236]), .D(n31), .Y(n466) );
  NAND2X1 U372 ( .A(n467), .B(n466), .Y(row[44]) );
  AOI22X1 U374 ( .A(regg[45]), .B(n3), .C(regg[109]), .D(n8), .Y(n472) );
  AOI22X1 U376 ( .A(regg[173]), .B(n41), .C(regg[237]), .D(n30), .Y(n471) );
  NAND2X1 U378 ( .A(n472), .B(n471), .Y(row[45]) );
  AOI22X1 U380 ( .A(regg[46]), .B(n2), .C(regg[110]), .D(n34), .Y(n474) );
  AOI22X1 U382 ( .A(regg[174]), .B(n43), .C(regg[238]), .D(n30), .Y(n473) );
  NAND2X1 U384 ( .A(n474), .B(n473), .Y(row[46]) );
  AOI22X1 U386 ( .A(regg[47]), .B(n3), .C(regg[111]), .D(n7), .Y(n476) );
  AOI22X1 U388 ( .A(regg[175]), .B(n45), .C(regg[239]), .D(n30), .Y(n475) );
  NAND2X1 U391 ( .A(n476), .B(n475), .Y(row[47]) );
  AOI22X1 U393 ( .A(regg[48]), .B(n14), .C(regg[112]), .D(n514), .Y(n478) );
  AOI22X1 U396 ( .A(regg[176]), .B(n32), .C(regg[240]), .D(n515), .Y(n477) );
  NAND2X1 U397 ( .A(n478), .B(n477), .Y(row[48]) );
  NAND2X1 U399 ( .A(regg[113]), .B(n514), .Y(n481) );
  NAND2X1 U401 ( .A(regg[241]), .B(n515), .Y(n480) );
  AOI22X1 U403 ( .A(regg[49]), .B(n14), .C(n32), .D(regg[177]), .Y(n479) );
  NAND3X1 U405 ( .A(n480), .B(n481), .C(n479), .Y(row[49]) );
  AOI22X1 U407 ( .A(n4), .B(regg[50]), .C(regg[114]), .D(n36), .Y(n483) );
  AOI22X1 U409 ( .A(n519), .B(regg[178]), .C(regg[242]), .D(n19), .Y(n482) );
  NAND2X1 U411 ( .A(n483), .B(n482), .Y(row[50]) );
  AOI22X1 U413 ( .A(regg[51]), .B(n37), .C(regg[115]), .D(n5), .Y(n488) );
  AOI22X1 U415 ( .A(regg[179]), .B(n44), .C(regg[243]), .D(n38), .Y(n487) );
  NAND2X1 U417 ( .A(n488), .B(n487), .Y(row[51]) );
  AOI22X1 U419 ( .A(regg[52]), .B(n12), .C(regg[116]), .D(n33), .Y(n490) );
  AOI22X1 U421 ( .A(regg[180]), .B(n44), .C(regg[244]), .D(n20), .Y(n489) );
  NAND2X1 U424 ( .A(n490), .B(n489), .Y(row[52]) );
  AOI22X1 U426 ( .A(regg[53]), .B(n12), .C(regg[117]), .D(n7), .Y(n492) );
  AOI22X1 U429 ( .A(regg[181]), .B(n45), .C(regg[245]), .D(n26), .Y(n491) );
  NAND2X1 U430 ( .A(n492), .B(n491), .Y(row[53]) );
  AOI22X1 U432 ( .A(regg[54]), .B(n9), .C(regg[118]), .D(n33), .Y(n494) );
  AOI22X1 U434 ( .A(regg[182]), .B(n41), .C(regg[246]), .D(n25), .Y(n493) );
  NAND2X1 U436 ( .A(n494), .B(n493), .Y(row[54]) );
  AOI22X1 U438 ( .A(regg[55]), .B(n37), .C(regg[119]), .D(n33), .Y(n496) );
  AOI22X1 U440 ( .A(regg[183]), .B(n43), .C(regg[247]), .D(n26), .Y(n495) );
  NAND2X1 U442 ( .A(n496), .B(n495), .Y(row[55]) );
  AOI22X1 U444 ( .A(regg[56]), .B(n9), .C(regg[120]), .D(n33), .Y(n498) );
  AOI22X1 U446 ( .A(regg[184]), .B(n43), .C(regg[248]), .D(n28), .Y(n497) );
  NAND2X1 U448 ( .A(n498), .B(n497), .Y(row[56]) );
  AOI22X1 U450 ( .A(regg[57]), .B(n37), .C(regg[121]), .D(n7), .Y(n503) );
  AOI22X1 U452 ( .A(regg[185]), .B(n45), .C(regg[249]), .D(n28), .Y(n499) );
  NAND2X1 U454 ( .A(n503), .B(n499), .Y(row[57]) );
  AOI22X1 U457 ( .A(regg[58]), .B(n9), .C(regg[122]), .D(n33), .Y(n505) );
  AOI22X1 U459 ( .A(regg[186]), .B(n41), .C(regg[250]), .D(n29), .Y(n504) );
  NAND2X1 U462 ( .A(n505), .B(n504), .Y(row[58]) );
  AOI22X1 U463 ( .A(regg[59]), .B(n2), .C(regg[123]), .D(n7), .Y(n507) );
  AOI22X1 U465 ( .A(regg[187]), .B(n45), .C(regg[251]), .D(n28), .Y(n506) );
  NAND2X1 U467 ( .A(n507), .B(n506), .Y(row[59]) );
  AOI22X1 U469 ( .A(regg[60]), .B(n9), .C(regg[124]), .D(n33), .Y(n509) );
  AOI22X1 U471 ( .A(regg[188]), .B(n45), .C(regg[252]), .D(n30), .Y(n508) );
  NAND2X1 U473 ( .A(n509), .B(n508), .Y(row[60]) );
  AOI22X1 U475 ( .A(regg[61]), .B(n2), .C(regg[125]), .D(n34), .Y(n511) );
  AOI22X1 U477 ( .A(regg[189]), .B(n43), .C(regg[253]), .D(n30), .Y(n510) );
  NAND2X1 U479 ( .A(n511), .B(n510), .Y(row[61]) );
  AOI22X1 U481 ( .A(regg[62]), .B(n2), .C(regg[126]), .D(n33), .Y(n513) );
  AOI22X1 U483 ( .A(regg[190]), .B(n41), .C(regg[254]), .D(n30), .Y(n512) );
  NAND2X1 U485 ( .A(n513), .B(n512), .Y(row[62]) );
  AOI22X1 U487 ( .A(regg[63]), .B(n9), .C(regg[127]), .D(n33), .Y(n521) );
  AOI22X1 U490 ( .A(regg[191]), .B(n45), .C(regg[255]), .D(n30), .Y(n520) );
  NAND2X1 U492 ( .A(n521), .B(n520), .Y(row[63]) );
  INVX2 U495 ( .A(n134), .Y(n522) );
  INVX2 U496 ( .A(n136), .Y(n523) );
  INVX2 U498 ( .A(n137), .Y(n524) );
  INVX2 U500 ( .A(n138), .Y(n525) );
  INVX2 U502 ( .A(n139), .Y(n526) );
  INVX2 U504 ( .A(n140), .Y(n527) );
  INVX2 U506 ( .A(n141), .Y(n528) );
  INVX2 U508 ( .A(n142), .Y(n529) );
  INVX2 U510 ( .A(n143), .Y(n530) );
  INVX2 U512 ( .A(n144), .Y(n531) );
  INVX2 U514 ( .A(n145), .Y(n535) );
  INVX2 U516 ( .A(n146), .Y(n536) );
  INVX2 U518 ( .A(n147), .Y(n537) );
  INVX2 U520 ( .A(n152), .Y(n538) );
  INVX2 U523 ( .A(n153), .Y(n539) );
  INVX2 U525 ( .A(n154), .Y(n540) );
  INVX2 U528 ( .A(n155), .Y(n541) );
  INVX2 U529 ( .A(n156), .Y(n542) );
  INVX2 U531 ( .A(n157), .Y(n543) );
  INVX2 U533 ( .A(n158), .Y(n544) );
  INVX2 U535 ( .A(n159), .Y(n545) );
  INVX2 U537 ( .A(n160), .Y(n546) );
  INVX2 U539 ( .A(n161), .Y(n547) );
  INVX2 U541 ( .A(n162), .Y(n551) );
  INVX2 U543 ( .A(n163), .Y(n552) );
  INVX2 U545 ( .A(n164), .Y(n553) );
  INVX2 U547 ( .A(n169), .Y(n554) );
  INVX2 U549 ( .A(n170), .Y(n555) );
  INVX2 U551 ( .A(n171), .Y(n556) );
  INVX2 U553 ( .A(n172), .Y(n557) );
  INVX2 U556 ( .A(n173), .Y(n558) );
  INVX2 U558 ( .A(n174), .Y(n559) );
  INVX2 U561 ( .A(n175), .Y(n560) );
  INVX2 U562 ( .A(n176), .Y(n561) );
  INVX2 U564 ( .A(n177), .Y(n562) );
  INVX2 U566 ( .A(n178), .Y(n563) );
  INVX2 U568 ( .A(n179), .Y(n567) );
  INVX2 U570 ( .A(n180), .Y(n568) );
  INVX2 U572 ( .A(n181), .Y(n569) );
  INVX2 U574 ( .A(n186), .Y(n570) );
  INVX2 U576 ( .A(n187), .Y(n571) );
  INVX2 U578 ( .A(n188), .Y(n572) );
  INVX2 U580 ( .A(n189), .Y(n573) );
  INVX2 U582 ( .A(n190), .Y(n574) );
  INVX2 U584 ( .A(n191), .Y(n575) );
  INVX2 U586 ( .A(n192), .Y(n576) );
  INVX2 U589 ( .A(n193), .Y(n577) );
  INVX2 U591 ( .A(n194), .Y(n578) );
  INVX2 U594 ( .A(n195), .Y(n579) );
  INVX2 U595 ( .A(n196), .Y(n583) );
  INVX2 U597 ( .A(n197), .Y(n584) );
  INVX2 U599 ( .A(n198), .Y(n585) );
  INVX2 U601 ( .A(n203), .Y(n586) );
  INVX2 U603 ( .A(n204), .Y(n587) );
  INVX2 U605 ( .A(n205), .Y(n588) );
  INVX2 U607 ( .A(n206), .Y(n589) );
  INVX2 U609 ( .A(n207), .Y(n590) );
  INVX2 U611 ( .A(n208), .Y(n591) );
  INVX2 U613 ( .A(n209), .Y(n592) );
  INVX2 U615 ( .A(n210), .Y(n593) );
  INVX2 U617 ( .A(n211), .Y(n594) );
  INVX2 U619 ( .A(n212), .Y(n595) );
  INVX2 U622 ( .A(n213), .Y(n599) );
  INVX2 U624 ( .A(n214), .Y(n600) );
  INVX2 U627 ( .A(n215), .Y(n601) );
  INVX2 U628 ( .A(n220), .Y(n602) );
  INVX2 U630 ( .A(n221), .Y(n603) );
  INVX2 U632 ( .A(n222), .Y(n604) );
  INVX2 U634 ( .A(n223), .Y(n605) );
  INVX2 U636 ( .A(n224), .Y(n606) );
  INVX2 U638 ( .A(n225), .Y(n607) );
  INVX2 U640 ( .A(n226), .Y(n608) );
  INVX2 U642 ( .A(n227), .Y(n609) );
  INVX2 U644 ( .A(n228), .Y(n610) );
  INVX2 U646 ( .A(n229), .Y(n611) );
  INVX2 U648 ( .A(n230), .Y(n615) );
  INVX2 U650 ( .A(n231), .Y(n616) );
  INVX2 U652 ( .A(n232), .Y(n617) );
  INVX2 U655 ( .A(n237), .Y(n618) );
  INVX2 U657 ( .A(n238), .Y(n619) );
  INVX2 U660 ( .A(n239), .Y(n620) );
  INVX2 U661 ( .A(n240), .Y(n621) );
  INVX2 U663 ( .A(n241), .Y(n622) );
  INVX2 U665 ( .A(n242), .Y(n623) );
  INVX2 U667 ( .A(n243), .Y(n624) );
  INVX2 U669 ( .A(n244), .Y(n625) );
  INVX2 U671 ( .A(n245), .Y(n626) );
  INVX2 U673 ( .A(n246), .Y(n627) );
  INVX2 U675 ( .A(n247), .Y(n631) );
  INVX2 U677 ( .A(n248), .Y(n632) );
  INVX2 U679 ( .A(n249), .Y(n633) );
  INVX2 U681 ( .A(n254), .Y(n634) );
  INVX2 U683 ( .A(n255), .Y(n635) );
  INVX2 U685 ( .A(n256), .Y(n636) );
  INVX2 U688 ( .A(n257), .Y(n637) );
  INVX2 U690 ( .A(n258), .Y(n638) );
  INVX2 U693 ( .A(n259), .Y(n639) );
  INVX2 U694 ( .A(n260), .Y(n640) );
  INVX2 U696 ( .A(n261), .Y(n641) );
  INVX2 U698 ( .A(n262), .Y(n642) );
  INVX2 U700 ( .A(n263), .Y(n643) );
  INVX2 U702 ( .A(n264), .Y(n647) );
  INVX2 U704 ( .A(n265), .Y(n648) );
  INVX2 U706 ( .A(n266), .Y(n649) );
  INVX2 U708 ( .A(n271), .Y(n650) );
  INVX2 U710 ( .A(n272), .Y(n651) );
  INVX2 U712 ( .A(n273), .Y(n652) );
  INVX2 U714 ( .A(n274), .Y(n653) );
  INVX2 U716 ( .A(n275), .Y(n654) );
  INVX2 U718 ( .A(n276), .Y(n655) );
  INVX2 U721 ( .A(n277), .Y(n656) );
  INVX2 U723 ( .A(n278), .Y(n657) );
  INVX2 U724 ( .A(n279), .Y(n658) );
  INVX2 U727 ( .A(n280), .Y(n659) );
  INVX2 U728 ( .A(n281), .Y(n663) );
  INVX2 U729 ( .A(n282), .Y(n664) );
  INVX2 U730 ( .A(n283), .Y(n665) );
  INVX2 U731 ( .A(n288), .Y(n666) );
  INVX2 U732 ( .A(n289), .Y(n667) );
  INVX2 U733 ( .A(n290), .Y(n668) );
  INVX2 U734 ( .A(n291), .Y(n669) );
  INVX2 U735 ( .A(n292), .Y(n670) );
  INVX2 U736 ( .A(n293), .Y(n671) );
  INVX2 U737 ( .A(n294), .Y(n672) );
  INVX2 U738 ( .A(n295), .Y(n673) );
  INVX2 U739 ( .A(n296), .Y(n674) );
  INVX2 U740 ( .A(n297), .Y(n675) );
  INVX2 U741 ( .A(n298), .Y(n676) );
  INVX2 U742 ( .A(n299), .Y(n677) );
  INVX2 U743 ( .A(n300), .Y(n678) );
  INVX2 U744 ( .A(n305), .Y(n679) );
  INVX2 U745 ( .A(n306), .Y(n680) );
  INVX2 U746 ( .A(n307), .Y(n681) );
  INVX2 U747 ( .A(n308), .Y(n682) );
  INVX2 U748 ( .A(n309), .Y(n683) );
  INVX2 U749 ( .A(n310), .Y(n684) );
  INVX2 U750 ( .A(n311), .Y(n685) );
  INVX2 U751 ( .A(n312), .Y(n686) );
  INVX2 U752 ( .A(n313), .Y(n687) );
  INVX2 U753 ( .A(n314), .Y(n688) );
  INVX2 U754 ( .A(n315), .Y(n689) );
  INVX2 U755 ( .A(n316), .Y(n690) );
  INVX2 U756 ( .A(n317), .Y(n691) );
  INVX2 U757 ( .A(n322), .Y(n692) );
  INVX2 U758 ( .A(n323), .Y(n693) );
  INVX2 U759 ( .A(n324), .Y(n694) );
  INVX2 U760 ( .A(n325), .Y(n695) );
  INVX2 U761 ( .A(n326), .Y(n696) );
  INVX2 U762 ( .A(n327), .Y(n697) );
  INVX2 U763 ( .A(n328), .Y(n698) );
  INVX2 U764 ( .A(n329), .Y(n699) );
  INVX2 U765 ( .A(n330), .Y(n700) );
  INVX2 U766 ( .A(n331), .Y(n701) );
  INVX2 U767 ( .A(n332), .Y(n702) );
  INVX2 U768 ( .A(n333), .Y(n703) );
  INVX2 U769 ( .A(n334), .Y(n704) );
  INVX2 U770 ( .A(n339), .Y(n705) );
  INVX2 U771 ( .A(n340), .Y(n706) );
  INVX2 U772 ( .A(n341), .Y(n707) );
  INVX2 U773 ( .A(n342), .Y(n708) );
  INVX2 U774 ( .A(n343), .Y(n709) );
  INVX2 U775 ( .A(n344), .Y(n710) );
  INVX2 U776 ( .A(n345), .Y(n711) );
  INVX2 U777 ( .A(n346), .Y(n712) );
  INVX2 U778 ( .A(n347), .Y(n713) );
  INVX2 U779 ( .A(n348), .Y(n714) );
  INVX2 U780 ( .A(n349), .Y(n715) );
  INVX2 U781 ( .A(n350), .Y(n716) );
  INVX2 U782 ( .A(n351), .Y(n717) );
  INVX2 U783 ( .A(n356), .Y(n718) );
  INVX2 U784 ( .A(n357), .Y(n719) );
  INVX2 U785 ( .A(n358), .Y(n720) );
  INVX2 U786 ( .A(n359), .Y(n721) );
  INVX2 U787 ( .A(n360), .Y(n722) );
  INVX2 U788 ( .A(n361), .Y(n723) );
  INVX2 U789 ( .A(n362), .Y(n724) );
  INVX2 U790 ( .A(n363), .Y(n725) );
  INVX2 U791 ( .A(n364), .Y(n726) );
  INVX2 U792 ( .A(n365), .Y(n727) );
  INVX2 U793 ( .A(n366), .Y(n728) );
  INVX2 U794 ( .A(n367), .Y(n729) );
  INVX2 U795 ( .A(n368), .Y(n730) );
  INVX2 U796 ( .A(n373), .Y(n731) );
  INVX2 U797 ( .A(n374), .Y(n732) );
  INVX2 U798 ( .A(n375), .Y(n733) );
  INVX2 U799 ( .A(n376), .Y(n734) );
  INVX2 U800 ( .A(n377), .Y(n735) );
  INVX2 U801 ( .A(n378), .Y(n736) );
  INVX2 U802 ( .A(n379), .Y(n737) );
  INVX2 U803 ( .A(n380), .Y(n738) );
  INVX2 U804 ( .A(n381), .Y(n739) );
  INVX2 U805 ( .A(n382), .Y(n740) );
  INVX2 U806 ( .A(n383), .Y(n741) );
  INVX2 U807 ( .A(n384), .Y(n742) );
  INVX2 U808 ( .A(n385), .Y(n743) );
  INVX2 U809 ( .A(n390), .Y(n744) );
  INVX2 U810 ( .A(n391), .Y(n745) );
  INVX2 U811 ( .A(n392), .Y(n746) );
  INVX2 U812 ( .A(n393), .Y(n747) );
  INVX2 U813 ( .A(n394), .Y(n748) );
  INVX2 U814 ( .A(n395), .Y(n749) );
  INVX2 U815 ( .A(n396), .Y(n750) );
  INVX2 U816 ( .A(n397), .Y(n751) );
  INVX2 U817 ( .A(n398), .Y(n752) );
  INVX2 U818 ( .A(n399), .Y(n753) );
  INVX2 U819 ( .A(n400), .Y(n754) );
  INVX2 U820 ( .A(n401), .Y(n755) );
  INVX2 U821 ( .A(n402), .Y(n756) );
  INVX2 U822 ( .A(regg[15]), .Y(n757) );
  INVX2 U823 ( .A(regg[31]), .Y(n758) );
  INVX2 U824 ( .A(regg[47]), .Y(n759) );
  INVX2 U825 ( .A(regg[14]), .Y(n760) );
  INVX2 U826 ( .A(regg[30]), .Y(n761) );
  INVX2 U827 ( .A(regg[46]), .Y(n762) );
  INVX2 U828 ( .A(regg[13]), .Y(n763) );
  INVX2 U829 ( .A(regg[29]), .Y(n764) );
  INVX2 U830 ( .A(regg[45]), .Y(n765) );
  INVX2 U831 ( .A(regg[12]), .Y(n766) );
  INVX2 U832 ( .A(regg[28]), .Y(n767) );
  INVX2 U833 ( .A(regg[44]), .Y(n768) );
  INVX2 U834 ( .A(regg[11]), .Y(n769) );
  INVX2 U835 ( .A(regg[27]), .Y(n770) );
  INVX2 U836 ( .A(regg[43]), .Y(n771) );
  INVX2 U837 ( .A(regg[10]), .Y(n772) );
  INVX2 U838 ( .A(regg[26]), .Y(n773) );
  INVX2 U839 ( .A(regg[42]), .Y(n774) );
  INVX2 U840 ( .A(regg[9]), .Y(n775) );
  INVX2 U841 ( .A(regg[25]), .Y(n776) );
  INVX2 U842 ( .A(regg[41]), .Y(n777) );
  INVX2 U843 ( .A(regg[8]), .Y(n778) );
  INVX2 U844 ( .A(regg[24]), .Y(n779) );
  INVX2 U845 ( .A(regg[40]), .Y(n780) );
  INVX2 U846 ( .A(regg[7]), .Y(n781) );
  INVX2 U847 ( .A(regg[23]), .Y(n782) );
  INVX2 U848 ( .A(regg[39]), .Y(n783) );
  INVX2 U849 ( .A(regg[6]), .Y(n784) );
  INVX2 U850 ( .A(regg[22]), .Y(n785) );
  INVX2 U851 ( .A(regg[38]), .Y(n786) );
  INVX2 U852 ( .A(regg[5]), .Y(n787) );
  INVX2 U853 ( .A(regg[21]), .Y(n788) );
  INVX2 U854 ( .A(regg[37]), .Y(n789) );
  INVX2 U855 ( .A(regg[4]), .Y(n790) );
  INVX2 U856 ( .A(regg[20]), .Y(n791) );
  INVX2 U857 ( .A(regg[36]), .Y(n792) );
  INVX2 U858 ( .A(regg[3]), .Y(n793) );
  INVX2 U859 ( .A(regg[19]), .Y(n794) );
  INVX2 U860 ( .A(regg[35]), .Y(n795) );
  INVX2 U861 ( .A(regg[2]), .Y(n796) );
  INVX2 U862 ( .A(regg[18]), .Y(n797) );
  INVX2 U863 ( .A(regg[34]), .Y(n798) );
  INVX2 U864 ( .A(regg[1]), .Y(n799) );
  INVX2 U865 ( .A(regg[17]), .Y(n800) );
  INVX2 U866 ( .A(regg[33]), .Y(n801) );
  INVX2 U867 ( .A(regg[0]), .Y(n802) );
  INVX2 U868 ( .A(regg[16]), .Y(n803) );
  INVX2 U869 ( .A(regg[32]), .Y(n804) );
endmodule


module coordinate_buffer ( strb_cor, databus_out, clk, sel, point );
  input [15:0] databus_out;
  output [47:0] point;
  input strb_cor, clk, sel;
  wire   n8, n15, n22, n29, n36, n43, n50, n57, n64, n71, n78, n85, n92, n99,
         n106, n113, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n1, n2,
         n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n16, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n30, n31, n32, n33, n34, n35,
         n37, n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n49, n51, n52,
         n53, n54, n55, n56, n58, n59, n60, n61, n62, n63, n65, n66, n67, n68,
         n69, n70, n72, n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84,
         n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97, n98, n100,
         n101, n102, n103, n104, n105, n107, n108, n109, n110, n111, n112,
         n114, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244;
  wire   [95:0] regg;
  tri   [15:0] databus_out;

  DFFPOSX1 \regg_reg[15]  ( .D(n210), .CLK(clk), .Q(regg[15]) );
  DFFPOSX1 \regg_reg[31]  ( .D(n209), .CLK(clk), .Q(regg[31]) );
  DFFPOSX1 \regg_reg[47]  ( .D(n208), .CLK(clk), .Q(regg[47]) );
  DFFPOSX1 \regg_reg[63]  ( .D(n207), .CLK(clk), .Q(regg[63]) );
  DFFPOSX1 \regg_reg[79]  ( .D(n206), .CLK(clk), .Q(regg[79]) );
  DFFPOSX1 \regg_reg[95]  ( .D(n205), .CLK(clk), .Q(regg[95]) );
  DFFPOSX1 \regg_reg[14]  ( .D(n204), .CLK(clk), .Q(regg[14]) );
  DFFPOSX1 \regg_reg[30]  ( .D(n203), .CLK(clk), .Q(regg[30]) );
  DFFPOSX1 \regg_reg[46]  ( .D(n202), .CLK(clk), .Q(regg[46]) );
  DFFPOSX1 \regg_reg[62]  ( .D(n201), .CLK(clk), .Q(regg[62]) );
  DFFPOSX1 \regg_reg[78]  ( .D(n200), .CLK(clk), .Q(regg[78]) );
  DFFPOSX1 \regg_reg[94]  ( .D(n199), .CLK(clk), .Q(regg[94]) );
  DFFPOSX1 \regg_reg[13]  ( .D(n198), .CLK(clk), .Q(regg[13]) );
  DFFPOSX1 \regg_reg[29]  ( .D(n197), .CLK(clk), .Q(regg[29]) );
  DFFPOSX1 \regg_reg[45]  ( .D(n196), .CLK(clk), .Q(regg[45]) );
  DFFPOSX1 \regg_reg[61]  ( .D(n195), .CLK(clk), .Q(regg[61]) );
  DFFPOSX1 \regg_reg[77]  ( .D(n194), .CLK(clk), .Q(regg[77]) );
  DFFPOSX1 \regg_reg[93]  ( .D(n193), .CLK(clk), .Q(regg[93]) );
  DFFPOSX1 \regg_reg[12]  ( .D(n192), .CLK(clk), .Q(regg[12]) );
  DFFPOSX1 \regg_reg[28]  ( .D(n191), .CLK(clk), .Q(regg[28]) );
  DFFPOSX1 \regg_reg[44]  ( .D(n190), .CLK(clk), .Q(regg[44]) );
  DFFPOSX1 \regg_reg[60]  ( .D(n189), .CLK(clk), .Q(regg[60]) );
  DFFPOSX1 \regg_reg[76]  ( .D(n188), .CLK(clk), .Q(regg[76]) );
  DFFPOSX1 \regg_reg[92]  ( .D(n187), .CLK(clk), .Q(regg[92]) );
  DFFPOSX1 \regg_reg[11]  ( .D(n186), .CLK(clk), .Q(regg[11]) );
  DFFPOSX1 \regg_reg[27]  ( .D(n185), .CLK(clk), .Q(regg[27]) );
  DFFPOSX1 \regg_reg[43]  ( .D(n184), .CLK(clk), .Q(regg[43]) );
  DFFPOSX1 \regg_reg[59]  ( .D(n183), .CLK(clk), .Q(regg[59]) );
  DFFPOSX1 \regg_reg[75]  ( .D(n182), .CLK(clk), .Q(regg[75]) );
  DFFPOSX1 \regg_reg[91]  ( .D(n181), .CLK(clk), .Q(regg[91]) );
  DFFPOSX1 \regg_reg[10]  ( .D(n180), .CLK(clk), .Q(regg[10]) );
  DFFPOSX1 \regg_reg[26]  ( .D(n179), .CLK(clk), .Q(regg[26]) );
  DFFPOSX1 \regg_reg[42]  ( .D(n178), .CLK(clk), .Q(regg[42]) );
  DFFPOSX1 \regg_reg[58]  ( .D(n177), .CLK(clk), .Q(regg[58]) );
  DFFPOSX1 \regg_reg[74]  ( .D(n176), .CLK(clk), .Q(regg[74]) );
  DFFPOSX1 \regg_reg[90]  ( .D(n175), .CLK(clk), .Q(regg[90]) );
  DFFPOSX1 \regg_reg[9]  ( .D(n174), .CLK(clk), .Q(regg[9]) );
  DFFPOSX1 \regg_reg[25]  ( .D(n173), .CLK(clk), .Q(regg[25]) );
  DFFPOSX1 \regg_reg[41]  ( .D(n172), .CLK(clk), .Q(regg[41]) );
  DFFPOSX1 \regg_reg[57]  ( .D(n171), .CLK(clk), .Q(regg[57]) );
  DFFPOSX1 \regg_reg[73]  ( .D(n170), .CLK(clk), .Q(regg[73]) );
  DFFPOSX1 \regg_reg[89]  ( .D(n169), .CLK(clk), .Q(regg[89]) );
  DFFPOSX1 \regg_reg[8]  ( .D(n168), .CLK(clk), .Q(regg[8]) );
  DFFPOSX1 \regg_reg[24]  ( .D(n167), .CLK(clk), .Q(regg[24]) );
  DFFPOSX1 \regg_reg[40]  ( .D(n166), .CLK(clk), .Q(regg[40]) );
  DFFPOSX1 \regg_reg[56]  ( .D(n165), .CLK(clk), .Q(regg[56]) );
  DFFPOSX1 \regg_reg[72]  ( .D(n164), .CLK(clk), .Q(regg[72]) );
  DFFPOSX1 \regg_reg[88]  ( .D(n163), .CLK(clk), .Q(regg[88]) );
  DFFPOSX1 \regg_reg[7]  ( .D(n162), .CLK(clk), .Q(regg[7]) );
  DFFPOSX1 \regg_reg[23]  ( .D(n161), .CLK(clk), .Q(regg[23]) );
  DFFPOSX1 \regg_reg[39]  ( .D(n160), .CLK(clk), .Q(regg[39]) );
  DFFPOSX1 \regg_reg[55]  ( .D(n159), .CLK(clk), .Q(regg[55]) );
  DFFPOSX1 \regg_reg[71]  ( .D(n158), .CLK(clk), .Q(regg[71]) );
  DFFPOSX1 \regg_reg[87]  ( .D(n157), .CLK(clk), .Q(regg[87]) );
  DFFPOSX1 \regg_reg[6]  ( .D(n156), .CLK(clk), .Q(regg[6]) );
  DFFPOSX1 \regg_reg[22]  ( .D(n155), .CLK(clk), .Q(regg[22]) );
  DFFPOSX1 \regg_reg[38]  ( .D(n154), .CLK(clk), .Q(regg[38]) );
  DFFPOSX1 \regg_reg[54]  ( .D(n153), .CLK(clk), .Q(regg[54]) );
  DFFPOSX1 \regg_reg[70]  ( .D(n152), .CLK(clk), .Q(regg[70]) );
  DFFPOSX1 \regg_reg[86]  ( .D(n151), .CLK(clk), .Q(regg[86]) );
  DFFPOSX1 \regg_reg[5]  ( .D(n150), .CLK(clk), .Q(regg[5]) );
  DFFPOSX1 \regg_reg[21]  ( .D(n149), .CLK(clk), .Q(regg[21]) );
  DFFPOSX1 \regg_reg[37]  ( .D(n148), .CLK(clk), .Q(regg[37]) );
  DFFPOSX1 \regg_reg[53]  ( .D(n147), .CLK(clk), .Q(regg[53]) );
  DFFPOSX1 \regg_reg[69]  ( .D(n146), .CLK(clk), .Q(regg[69]) );
  DFFPOSX1 \regg_reg[85]  ( .D(n145), .CLK(clk), .Q(regg[85]) );
  DFFPOSX1 \regg_reg[4]  ( .D(n144), .CLK(clk), .Q(regg[4]) );
  DFFPOSX1 \regg_reg[20]  ( .D(n143), .CLK(clk), .Q(regg[20]) );
  DFFPOSX1 \regg_reg[36]  ( .D(n142), .CLK(clk), .Q(regg[36]) );
  DFFPOSX1 \regg_reg[52]  ( .D(n141), .CLK(clk), .Q(regg[52]) );
  DFFPOSX1 \regg_reg[68]  ( .D(n140), .CLK(clk), .Q(regg[68]) );
  DFFPOSX1 \regg_reg[84]  ( .D(n139), .CLK(clk), .Q(regg[84]) );
  DFFPOSX1 \regg_reg[3]  ( .D(n138), .CLK(clk), .Q(regg[3]) );
  DFFPOSX1 \regg_reg[19]  ( .D(n137), .CLK(clk), .Q(regg[19]) );
  DFFPOSX1 \regg_reg[35]  ( .D(n136), .CLK(clk), .Q(regg[35]) );
  DFFPOSX1 \regg_reg[51]  ( .D(n135), .CLK(clk), .Q(regg[51]) );
  DFFPOSX1 \regg_reg[67]  ( .D(n134), .CLK(clk), .Q(regg[67]) );
  DFFPOSX1 \regg_reg[83]  ( .D(n133), .CLK(clk), .Q(regg[83]) );
  DFFPOSX1 \regg_reg[2]  ( .D(n132), .CLK(clk), .Q(regg[2]) );
  DFFPOSX1 \regg_reg[18]  ( .D(n131), .CLK(clk), .Q(regg[18]) );
  DFFPOSX1 \regg_reg[34]  ( .D(n130), .CLK(clk), .Q(regg[34]) );
  DFFPOSX1 \regg_reg[50]  ( .D(n129), .CLK(clk), .Q(regg[50]) );
  DFFPOSX1 \regg_reg[66]  ( .D(n128), .CLK(clk), .Q(regg[66]) );
  DFFPOSX1 \regg_reg[82]  ( .D(n127), .CLK(clk), .Q(regg[82]) );
  DFFPOSX1 \regg_reg[1]  ( .D(n126), .CLK(clk), .Q(regg[1]) );
  DFFPOSX1 \regg_reg[17]  ( .D(n125), .CLK(clk), .Q(regg[17]) );
  DFFPOSX1 \regg_reg[33]  ( .D(n124), .CLK(clk), .Q(regg[33]) );
  DFFPOSX1 \regg_reg[49]  ( .D(n123), .CLK(clk), .Q(regg[49]) );
  DFFPOSX1 \regg_reg[65]  ( .D(n122), .CLK(clk), .Q(regg[65]) );
  DFFPOSX1 \regg_reg[81]  ( .D(n121), .CLK(clk), .Q(regg[81]) );
  DFFPOSX1 \regg_reg[0]  ( .D(n120), .CLK(clk), .Q(regg[0]) );
  DFFPOSX1 \regg_reg[16]  ( .D(n119), .CLK(clk), .Q(regg[16]) );
  DFFPOSX1 \regg_reg[32]  ( .D(n118), .CLK(clk), .Q(regg[32]) );
  DFFPOSX1 \regg_reg[48]  ( .D(n117), .CLK(clk), .Q(regg[48]) );
  DFFPOSX1 \regg_reg[64]  ( .D(n116), .CLK(clk), .Q(regg[64]) );
  DFFPOSX1 \regg_reg[80]  ( .D(n115), .CLK(clk), .Q(regg[80]) );
  NAND2X1 U8 ( .A(databus_out[0]), .B(n11), .Y(n8) );
  NAND2X1 U15 ( .A(databus_out[1]), .B(n13), .Y(n15) );
  NAND2X1 U22 ( .A(databus_out[2]), .B(n10), .Y(n22) );
  NAND2X1 U29 ( .A(databus_out[3]), .B(n12), .Y(n29) );
  NAND2X1 U36 ( .A(databus_out[4]), .B(n14), .Y(n36) );
  NAND2X1 U43 ( .A(databus_out[5]), .B(n11), .Y(n43) );
  NAND2X1 U50 ( .A(databus_out[6]), .B(n13), .Y(n50) );
  NAND2X1 U57 ( .A(databus_out[7]), .B(n11), .Y(n57) );
  NAND2X1 U64 ( .A(databus_out[8]), .B(n16), .Y(n64) );
  NAND2X1 U71 ( .A(databus_out[9]), .B(n13), .Y(n71) );
  NAND2X1 U78 ( .A(databus_out[10]), .B(n9), .Y(n78) );
  NAND2X1 U85 ( .A(databus_out[11]), .B(n9), .Y(n85) );
  NAND2X1 U92 ( .A(databus_out[12]), .B(n9), .Y(n92) );
  NAND2X1 U99 ( .A(databus_out[13]), .B(n10), .Y(n99) );
  NAND2X1 U106 ( .A(databus_out[14]), .B(n12), .Y(n106) );
  NAND2X1 U114 ( .A(databus_out[15]), .B(n9), .Y(n113) );
  INVX2 U2 ( .A(n4), .Y(n2) );
  INVX1 U3 ( .A(n40), .Y(n1) );
  BUFX4 U4 ( .A(sel), .Y(n3) );
  INVX2 U5 ( .A(sel), .Y(n40) );
  MUX2X1 U6 ( .B(n111), .A(n108), .S(n40), .Y(point[9]) );
  MUX2X1 U7 ( .B(n237), .A(n234), .S(n40), .Y(point[30]) );
  MUX2X1 U9 ( .B(n232), .A(n229), .S(n40), .Y(point[13]) );
  MUX2X1 U10 ( .B(n213), .A(n114), .S(n40), .Y(point[26]) );
  BUFX4 U11 ( .A(sel), .Y(n4) );
  MUX2X1 U12 ( .B(n62), .A(n59), .S(n2), .Y(point[2]) );
  INVX2 U13 ( .A(n25), .Y(n10) );
  INVX2 U14 ( .A(n19), .Y(n16) );
  INVX2 U16 ( .A(n20), .Y(n14) );
  INVX2 U17 ( .A(n21), .Y(n13) );
  INVX2 U18 ( .A(n24), .Y(n11) );
  INVX2 U19 ( .A(n23), .Y(n12) );
  INVX2 U20 ( .A(n26), .Y(n9) );
  BUFX2 U21 ( .A(n37), .Y(n19) );
  BUFX2 U23 ( .A(n37), .Y(n20) );
  BUFX2 U24 ( .A(n37), .Y(n21) );
  BUFX2 U25 ( .A(n37), .Y(n23) );
  BUFX2 U26 ( .A(n37), .Y(n24) );
  BUFX2 U27 ( .A(n37), .Y(n25) );
  BUFX2 U28 ( .A(n37), .Y(n26) );
  BUFX2 U30 ( .A(n37), .Y(n17) );
  BUFX2 U31 ( .A(n37), .Y(n18) );
  BUFX2 U32 ( .A(n17), .Y(n27) );
  BUFX2 U33 ( .A(n17), .Y(n28) );
  BUFX2 U34 ( .A(n17), .Y(n30) );
  BUFX2 U35 ( .A(n37), .Y(n31) );
  BUFX2 U37 ( .A(n37), .Y(n32) );
  BUFX2 U38 ( .A(n37), .Y(n33) );
  BUFX2 U39 ( .A(n37), .Y(n34) );
  BUFX2 U40 ( .A(n37), .Y(n35) );
  INVX2 U41 ( .A(strb_cor), .Y(n37) );
  INVX4 U42 ( .A(n6), .Y(point[31]) );
  INVX4 U44 ( .A(n7), .Y(point[15]) );
  INVX4 U45 ( .A(n5), .Y(point[47]) );
  MUX2X1 U46 ( .B(regg[95]), .A(regg[47]), .S(n38), .Y(n5) );
  INVX1 U47 ( .A(regg[95]), .Y(n239) );
  INVX1 U48 ( .A(regg[47]), .Y(n242) );
  INVX4 U49 ( .A(sel), .Y(n41) );
  MUX2X1 U51 ( .B(regg[31]), .A(regg[79]), .S(n2), .Y(n6) );
  INVX1 U52 ( .A(regg[31]), .Y(n243) );
  INVX1 U53 ( .A(regg[79]), .Y(n240) );
  MUX2X1 U54 ( .B(regg[15]), .A(regg[63]), .S(n40), .Y(n7) );
  INVX1 U55 ( .A(regg[15]), .Y(n244) );
  INVX1 U56 ( .A(regg[63]), .Y(n241) );
  INVX8 U58 ( .A(n41), .Y(n38) );
  INVX8 U59 ( .A(n41), .Y(n39) );
  INVX2 U60 ( .A(regg[48]), .Y(n45) );
  INVX2 U61 ( .A(regg[0]), .Y(n48) );
  MUX2X1 U62 ( .B(n45), .A(n48), .S(n38), .Y(point[0]) );
  INVX2 U63 ( .A(regg[49]), .Y(n52) );
  INVX2 U65 ( .A(regg[1]), .Y(n55) );
  MUX2X1 U66 ( .B(n52), .A(n55), .S(n38), .Y(point[1]) );
  INVX2 U67 ( .A(regg[50]), .Y(n59) );
  INVX2 U68 ( .A(regg[2]), .Y(n62) );
  INVX2 U69 ( .A(regg[51]), .Y(n66) );
  INVX2 U70 ( .A(regg[3]), .Y(n69) );
  MUX2X1 U72 ( .B(n66), .A(n69), .S(n38), .Y(point[3]) );
  INVX2 U73 ( .A(regg[52]), .Y(n73) );
  INVX2 U74 ( .A(regg[4]), .Y(n76) );
  MUX2X1 U75 ( .B(n73), .A(n76), .S(n38), .Y(point[4]) );
  INVX2 U76 ( .A(regg[53]), .Y(n80) );
  INVX2 U77 ( .A(regg[5]), .Y(n83) );
  MUX2X1 U79 ( .B(n80), .A(n83), .S(n38), .Y(point[5]) );
  INVX2 U80 ( .A(regg[54]), .Y(n87) );
  INVX2 U81 ( .A(regg[6]), .Y(n90) );
  MUX2X1 U82 ( .B(n87), .A(n90), .S(n38), .Y(point[6]) );
  INVX2 U83 ( .A(regg[55]), .Y(n94) );
  INVX2 U84 ( .A(regg[7]), .Y(n97) );
  MUX2X1 U86 ( .B(n94), .A(n97), .S(n38), .Y(point[7]) );
  INVX2 U87 ( .A(regg[56]), .Y(n101) );
  INVX2 U88 ( .A(regg[8]), .Y(n104) );
  MUX2X1 U89 ( .B(n101), .A(n104), .S(n39), .Y(point[8]) );
  INVX2 U90 ( .A(regg[57]), .Y(n108) );
  INVX2 U91 ( .A(regg[9]), .Y(n111) );
  INVX2 U93 ( .A(regg[58]), .Y(n211) );
  INVX2 U94 ( .A(regg[10]), .Y(n214) );
  MUX2X1 U95 ( .B(n211), .A(n214), .S(n38), .Y(point[10]) );
  INVX2 U96 ( .A(regg[59]), .Y(n217) );
  INVX2 U97 ( .A(regg[11]), .Y(n220) );
  MUX2X1 U98 ( .B(n217), .A(n220), .S(n4), .Y(point[11]) );
  INVX2 U100 ( .A(regg[60]), .Y(n223) );
  INVX2 U101 ( .A(regg[12]), .Y(n226) );
  MUX2X1 U102 ( .B(n223), .A(n226), .S(n3), .Y(point[12]) );
  INVX2 U103 ( .A(regg[61]), .Y(n229) );
  INVX2 U104 ( .A(regg[13]), .Y(n232) );
  INVX2 U105 ( .A(regg[62]), .Y(n235) );
  INVX2 U107 ( .A(regg[14]), .Y(n238) );
  MUX2X1 U108 ( .B(n235), .A(n238), .S(n39), .Y(point[14]) );
  INVX2 U109 ( .A(regg[64]), .Y(n44) );
  INVX2 U110 ( .A(regg[16]), .Y(n47) );
  MUX2X1 U111 ( .B(n44), .A(n47), .S(n38), .Y(point[16]) );
  INVX2 U112 ( .A(regg[65]), .Y(n51) );
  INVX2 U113 ( .A(regg[17]), .Y(n54) );
  MUX2X1 U115 ( .B(n51), .A(n54), .S(n38), .Y(point[17]) );
  INVX2 U116 ( .A(regg[66]), .Y(n58) );
  INVX2 U117 ( .A(regg[18]), .Y(n61) );
  MUX2X1 U118 ( .B(n58), .A(n61), .S(n38), .Y(point[18]) );
  INVX2 U119 ( .A(regg[67]), .Y(n65) );
  INVX2 U120 ( .A(regg[19]), .Y(n68) );
  MUX2X1 U121 ( .B(n65), .A(n68), .S(n38), .Y(point[19]) );
  INVX2 U122 ( .A(regg[68]), .Y(n72) );
  INVX2 U123 ( .A(regg[20]), .Y(n75) );
  MUX2X1 U124 ( .B(n72), .A(n75), .S(n39), .Y(point[20]) );
  INVX2 U125 ( .A(regg[69]), .Y(n79) );
  INVX2 U126 ( .A(regg[21]), .Y(n82) );
  MUX2X1 U127 ( .B(n79), .A(n82), .S(n39), .Y(point[21]) );
  INVX2 U128 ( .A(regg[70]), .Y(n86) );
  INVX2 U129 ( .A(regg[22]), .Y(n89) );
  MUX2X1 U130 ( .B(n86), .A(n89), .S(n39), .Y(point[22]) );
  INVX2 U131 ( .A(regg[71]), .Y(n93) );
  INVX2 U132 ( .A(regg[23]), .Y(n96) );
  MUX2X1 U133 ( .B(n93), .A(n96), .S(n38), .Y(point[23]) );
  INVX2 U134 ( .A(regg[72]), .Y(n100) );
  INVX2 U135 ( .A(regg[24]), .Y(n103) );
  MUX2X1 U136 ( .B(n100), .A(n103), .S(n3), .Y(point[24]) );
  INVX2 U137 ( .A(regg[73]), .Y(n107) );
  INVX2 U138 ( .A(regg[25]), .Y(n110) );
  MUX2X1 U139 ( .B(n107), .A(n110), .S(n4), .Y(point[25]) );
  INVX2 U140 ( .A(regg[74]), .Y(n114) );
  INVX2 U141 ( .A(regg[26]), .Y(n213) );
  INVX2 U142 ( .A(regg[75]), .Y(n216) );
  INVX2 U143 ( .A(regg[27]), .Y(n219) );
  MUX2X1 U144 ( .B(n216), .A(n219), .S(n39), .Y(point[27]) );
  INVX2 U145 ( .A(regg[76]), .Y(n222) );
  INVX2 U146 ( .A(regg[28]), .Y(n225) );
  MUX2X1 U147 ( .B(n222), .A(n225), .S(n4), .Y(point[28]) );
  INVX2 U148 ( .A(regg[77]), .Y(n228) );
  INVX2 U149 ( .A(regg[29]), .Y(n231) );
  MUX2X1 U150 ( .B(n228), .A(n231), .S(n39), .Y(point[29]) );
  INVX2 U151 ( .A(regg[78]), .Y(n234) );
  INVX2 U152 ( .A(regg[30]), .Y(n237) );
  INVX2 U153 ( .A(regg[80]), .Y(n42) );
  INVX2 U154 ( .A(regg[32]), .Y(n46) );
  MUX2X1 U155 ( .B(n42), .A(n46), .S(n38), .Y(point[32]) );
  INVX2 U156 ( .A(regg[81]), .Y(n49) );
  INVX2 U157 ( .A(regg[33]), .Y(n53) );
  MUX2X1 U158 ( .B(n49), .A(n53), .S(n38), .Y(point[33]) );
  INVX2 U159 ( .A(regg[82]), .Y(n56) );
  INVX2 U160 ( .A(regg[34]), .Y(n60) );
  MUX2X1 U161 ( .B(n56), .A(n60), .S(n38), .Y(point[34]) );
  INVX2 U162 ( .A(regg[83]), .Y(n63) );
  INVX2 U163 ( .A(regg[35]), .Y(n67) );
  MUX2X1 U164 ( .B(n63), .A(n67), .S(n38), .Y(point[35]) );
  INVX2 U165 ( .A(regg[84]), .Y(n70) );
  INVX2 U166 ( .A(regg[36]), .Y(n74) );
  MUX2X1 U167 ( .B(n70), .A(n74), .S(n39), .Y(point[36]) );
  INVX2 U168 ( .A(regg[85]), .Y(n77) );
  INVX2 U169 ( .A(regg[37]), .Y(n81) );
  MUX2X1 U170 ( .B(n77), .A(n81), .S(n38), .Y(point[37]) );
  INVX2 U171 ( .A(regg[86]), .Y(n84) );
  INVX2 U172 ( .A(regg[38]), .Y(n88) );
  MUX2X1 U173 ( .B(n84), .A(n88), .S(n3), .Y(point[38]) );
  INVX2 U174 ( .A(regg[87]), .Y(n91) );
  INVX2 U175 ( .A(regg[39]), .Y(n95) );
  MUX2X1 U176 ( .B(n91), .A(n95), .S(n3), .Y(point[39]) );
  INVX2 U177 ( .A(regg[88]), .Y(n98) );
  INVX2 U178 ( .A(regg[40]), .Y(n102) );
  MUX2X1 U179 ( .B(n98), .A(n102), .S(n3), .Y(point[40]) );
  INVX2 U180 ( .A(regg[89]), .Y(n105) );
  INVX2 U181 ( .A(regg[41]), .Y(n109) );
  MUX2X1 U182 ( .B(n105), .A(n109), .S(n3), .Y(point[41]) );
  INVX2 U183 ( .A(regg[90]), .Y(n112) );
  INVX2 U184 ( .A(regg[42]), .Y(n212) );
  MUX2X1 U185 ( .B(n112), .A(n212), .S(n39), .Y(point[42]) );
  INVX2 U186 ( .A(regg[91]), .Y(n215) );
  INVX2 U187 ( .A(regg[43]), .Y(n218) );
  MUX2X1 U188 ( .B(n215), .A(n218), .S(n4), .Y(point[43]) );
  INVX2 U189 ( .A(regg[92]), .Y(n221) );
  INVX2 U190 ( .A(regg[44]), .Y(n224) );
  MUX2X1 U191 ( .B(n221), .A(n224), .S(n1), .Y(point[44]) );
  INVX2 U192 ( .A(regg[93]), .Y(n227) );
  INVX2 U193 ( .A(regg[45]), .Y(n230) );
  MUX2X1 U194 ( .B(n227), .A(n230), .S(n39), .Y(point[45]) );
  INVX2 U195 ( .A(regg[94]), .Y(n233) );
  INVX2 U196 ( .A(regg[46]), .Y(n236) );
  MUX2X1 U197 ( .B(n233), .A(n236), .S(n38), .Y(point[46]) );
  OAI22X1 U198 ( .A(n42), .B(n13), .C(n17), .D(n44), .Y(n115) );
  OAI22X1 U199 ( .A(n44), .B(n12), .C(n17), .D(n45), .Y(n116) );
  OAI22X1 U200 ( .A(n45), .B(n10), .C(n17), .D(n46), .Y(n117) );
  OAI22X1 U201 ( .A(n46), .B(n13), .C(n18), .D(n47), .Y(n118) );
  OAI22X1 U202 ( .A(n47), .B(n11), .C(n18), .D(n48), .Y(n119) );
  OAI21X1 U203 ( .A(n48), .B(n9), .C(n8), .Y(n120) );
  OAI22X1 U204 ( .A(n49), .B(n16), .C(n18), .D(n51), .Y(n121) );
  OAI22X1 U205 ( .A(n51), .B(n14), .C(n19), .D(n52), .Y(n122) );
  OAI22X1 U206 ( .A(n52), .B(n16), .C(n19), .D(n53), .Y(n123) );
  OAI22X1 U207 ( .A(n53), .B(n16), .C(n19), .D(n54), .Y(n124) );
  OAI22X1 U208 ( .A(n54), .B(n16), .C(n20), .D(n55), .Y(n125) );
  OAI21X1 U209 ( .A(n55), .B(n9), .C(n15), .Y(n126) );
  OAI22X1 U210 ( .A(n56), .B(n16), .C(n20), .D(n58), .Y(n127) );
  OAI22X1 U211 ( .A(n58), .B(n16), .C(n20), .D(n59), .Y(n128) );
  OAI22X1 U212 ( .A(n59), .B(n16), .C(n21), .D(n60), .Y(n129) );
  OAI22X1 U213 ( .A(n60), .B(n16), .C(n21), .D(n61), .Y(n130) );
  OAI22X1 U214 ( .A(n61), .B(n16), .C(n21), .D(n62), .Y(n131) );
  OAI21X1 U215 ( .A(n62), .B(n9), .C(n22), .Y(n132) );
  OAI22X1 U216 ( .A(n63), .B(n16), .C(n23), .D(n65), .Y(n133) );
  OAI22X1 U217 ( .A(n65), .B(n16), .C(n23), .D(n66), .Y(n134) );
  OAI22X1 U218 ( .A(n66), .B(n16), .C(n23), .D(n67), .Y(n135) );
  OAI22X1 U219 ( .A(n67), .B(n16), .C(n24), .D(n68), .Y(n136) );
  OAI22X1 U220 ( .A(n68), .B(n16), .C(n24), .D(n69), .Y(n137) );
  OAI21X1 U221 ( .A(n69), .B(n9), .C(n29), .Y(n138) );
  OAI22X1 U222 ( .A(n70), .B(n14), .C(n24), .D(n72), .Y(n139) );
  OAI22X1 U223 ( .A(n72), .B(n14), .C(n25), .D(n73), .Y(n140) );
  OAI22X1 U224 ( .A(n73), .B(n14), .C(n25), .D(n74), .Y(n141) );
  OAI22X1 U225 ( .A(n74), .B(n14), .C(n25), .D(n75), .Y(n142) );
  OAI22X1 U226 ( .A(n75), .B(n14), .C(n26), .D(n76), .Y(n143) );
  OAI21X1 U227 ( .A(n76), .B(n10), .C(n36), .Y(n144) );
  OAI22X1 U228 ( .A(n77), .B(n14), .C(n26), .D(n79), .Y(n145) );
  OAI22X1 U229 ( .A(n79), .B(n14), .C(n26), .D(n80), .Y(n146) );
  OAI22X1 U230 ( .A(n80), .B(n14), .C(n27), .D(n81), .Y(n147) );
  OAI22X1 U231 ( .A(n81), .B(n14), .C(n27), .D(n82), .Y(n148) );
  OAI22X1 U232 ( .A(n82), .B(n14), .C(n27), .D(n83), .Y(n149) );
  OAI21X1 U233 ( .A(n83), .B(n9), .C(n43), .Y(n150) );
  OAI22X1 U234 ( .A(n84), .B(n14), .C(n27), .D(n86), .Y(n151) );
  OAI22X1 U235 ( .A(n86), .B(n14), .C(n27), .D(n87), .Y(n152) );
  OAI22X1 U236 ( .A(n87), .B(n14), .C(n27), .D(n88), .Y(n153) );
  OAI22X1 U237 ( .A(n88), .B(n13), .C(n27), .D(n89), .Y(n154) );
  OAI22X1 U238 ( .A(n89), .B(n13), .C(n28), .D(n90), .Y(n155) );
  OAI21X1 U239 ( .A(n90), .B(n9), .C(n50), .Y(n156) );
  OAI22X1 U240 ( .A(n91), .B(n13), .C(n28), .D(n93), .Y(n157) );
  OAI22X1 U241 ( .A(n93), .B(n13), .C(n28), .D(n94), .Y(n158) );
  OAI22X1 U242 ( .A(n94), .B(n13), .C(n28), .D(n95), .Y(n159) );
  OAI22X1 U243 ( .A(n95), .B(n13), .C(n28), .D(n96), .Y(n160) );
  OAI22X1 U244 ( .A(n96), .B(n13), .C(n28), .D(n97), .Y(n161) );
  OAI21X1 U245 ( .A(n97), .B(n9), .C(n57), .Y(n162) );
  OAI22X1 U246 ( .A(n98), .B(n13), .C(n28), .D(n100), .Y(n163) );
  OAI22X1 U247 ( .A(n100), .B(n13), .C(n30), .D(n101), .Y(n164) );
  OAI22X1 U248 ( .A(n101), .B(n13), .C(n30), .D(n102), .Y(n165) );
  OAI22X1 U249 ( .A(n102), .B(n13), .C(n30), .D(n103), .Y(n166) );
  OAI22X1 U250 ( .A(n103), .B(n13), .C(n30), .D(n104), .Y(n167) );
  OAI21X1 U251 ( .A(n104), .B(n10), .C(n64), .Y(n168) );
  OAI22X1 U252 ( .A(n105), .B(n12), .C(n30), .D(n107), .Y(n169) );
  OAI22X1 U253 ( .A(n107), .B(n12), .C(n30), .D(n108), .Y(n170) );
  OAI22X1 U254 ( .A(n108), .B(n12), .C(n30), .D(n109), .Y(n171) );
  OAI22X1 U255 ( .A(n109), .B(n12), .C(n31), .D(n110), .Y(n172) );
  OAI22X1 U256 ( .A(n110), .B(n12), .C(n31), .D(n111), .Y(n173) );
  OAI21X1 U257 ( .A(n111), .B(n9), .C(n71), .Y(n174) );
  OAI22X1 U258 ( .A(n112), .B(n12), .C(n31), .D(n114), .Y(n175) );
  OAI22X1 U259 ( .A(n114), .B(n12), .C(n31), .D(n211), .Y(n176) );
  OAI22X1 U260 ( .A(n211), .B(n12), .C(n31), .D(n212), .Y(n177) );
  OAI22X1 U261 ( .A(n212), .B(n12), .C(n31), .D(n213), .Y(n178) );
  OAI22X1 U262 ( .A(n213), .B(n12), .C(n31), .D(n214), .Y(n179) );
  OAI21X1 U263 ( .A(n214), .B(n10), .C(n78), .Y(n180) );
  OAI22X1 U264 ( .A(n215), .B(n11), .C(n32), .D(n216), .Y(n181) );
  OAI22X1 U265 ( .A(n216), .B(n11), .C(n32), .D(n217), .Y(n182) );
  OAI22X1 U266 ( .A(n217), .B(n11), .C(n32), .D(n218), .Y(n183) );
  OAI22X1 U267 ( .A(n218), .B(n12), .C(n32), .D(n219), .Y(n184) );
  OAI22X1 U268 ( .A(n219), .B(n11), .C(n32), .D(n220), .Y(n185) );
  OAI21X1 U269 ( .A(n220), .B(n10), .C(n85), .Y(n186) );
  OAI22X1 U270 ( .A(n221), .B(n12), .C(n32), .D(n222), .Y(n187) );
  OAI22X1 U271 ( .A(n222), .B(n11), .C(n32), .D(n223), .Y(n188) );
  OAI22X1 U272 ( .A(n223), .B(n11), .C(n33), .D(n224), .Y(n189) );
  OAI22X1 U273 ( .A(n224), .B(n11), .C(n33), .D(n225), .Y(n190) );
  OAI22X1 U274 ( .A(n225), .B(n11), .C(n33), .D(n226), .Y(n191) );
  OAI21X1 U275 ( .A(n226), .B(n9), .C(n92), .Y(n192) );
  OAI22X1 U276 ( .A(n227), .B(n11), .C(n33), .D(n228), .Y(n193) );
  OAI22X1 U277 ( .A(n228), .B(n11), .C(n33), .D(n229), .Y(n194) );
  OAI22X1 U278 ( .A(n229), .B(n11), .C(n33), .D(n230), .Y(n195) );
  OAI22X1 U279 ( .A(n230), .B(n10), .C(n33), .D(n231), .Y(n196) );
  OAI22X1 U280 ( .A(n231), .B(n11), .C(n34), .D(n232), .Y(n197) );
  OAI21X1 U281 ( .A(n232), .B(n9), .C(n99), .Y(n198) );
  OAI22X1 U282 ( .A(n233), .B(n10), .C(n34), .D(n234), .Y(n199) );
  OAI22X1 U283 ( .A(n234), .B(n10), .C(n34), .D(n235), .Y(n200) );
  OAI22X1 U284 ( .A(n235), .B(n10), .C(n34), .D(n236), .Y(n201) );
  OAI22X1 U285 ( .A(n236), .B(n10), .C(n34), .D(n237), .Y(n202) );
  OAI22X1 U286 ( .A(n237), .B(n10), .C(n34), .D(n238), .Y(n203) );
  OAI21X1 U287 ( .A(n238), .B(n9), .C(n106), .Y(n204) );
  OAI22X1 U288 ( .A(n239), .B(n10), .C(n34), .D(n240), .Y(n205) );
  OAI22X1 U289 ( .A(n240), .B(n10), .C(n35), .D(n241), .Y(n206) );
  OAI22X1 U290 ( .A(n241), .B(n11), .C(n35), .D(n242), .Y(n207) );
  OAI22X1 U291 ( .A(n242), .B(n10), .C(n35), .D(n243), .Y(n208) );
  OAI22X1 U292 ( .A(n243), .B(n12), .C(n35), .D(n244), .Y(n209) );
  OAI21X1 U293 ( .A(n244), .B(n9), .C(n113), .Y(n210) );
endmodule


module gpu_controller_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
endmodule


module gpu_controller ( databus, strb_in, clk, rst_n, gpu_done, ram_in_use, 
        rast_done, init_rast, rast_addr, rast_strb, rast_index, math_done, 
        init_math, strb_matrix, strb_cor, err, addr_out, re_out, we_out, 
        databus_out, opp );
  inout [15:0] databus;
  input [15:0] rast_addr;
  input [3:0] rast_index;
  output [14:0] addr_out;
  output [15:0] databus_out;
  output [15:0] opp;
  input strb_in, clk, rst_n, ram_in_use, rast_done, rast_strb, math_done, err;
  output gpu_done, init_rast, init_math, strb_matrix, strb_cor, re_out, we_out;
  wire   re, we, tem, tem2, nextre, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N314, N315,
         N316, N317, n1, n2, n3, n7, n8, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n48,
         n49, n51, n52, n53, n54, n59, n61, n63, n65, n67, n68, n69, n73, n74,
         n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n90,
         n91, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n104, n105,
         n107, n108, n109, n110, n111, n112, n114, n115, n116, n117, n119,
         n120, n122, n123, n124, n126, n127, n128, n129, n130, n132, n133,
         n134, n135, n137, n138, n140, n141, n142, n143, n144, n146, n147,
         n149, n150, n151, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n165, n166, n167, n169, n170, n171, n172, n173, n174,
         n176, n177, n178, n180, n182, n183, n184, n185, n186, n187, n189,
         n190, n193, n194, n195, n196, n197, n198, n199, n200, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n274, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n293, n294, n295, n296, n297, n298, n300, n312, n314,
         n324, n326, n328, n329, n330, n331, \add_213/carry[4] ,
         \add_213/carry[3] , \add_213/carry[2] , n4, n5, n6, n9, n10, n11, n12,
         n47, n50, n55, n56, n57, n58, n60, n62, n64, n66, n70, n71, n72, n76,
         n89, n92, n103, n106, n113, n118, n121, n125, n131, n136, n139, n145,
         n148, n152, n153, n164, n168, n175, n179, n181, n188, n191, n192,
         n201, n211, n212, n213, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n275, n292, n299, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n313,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n325, n327,
         n332, n333;
  wire   [3:0] state;
  wire   [15:0] addr;
  wire   [4:0] counter;
  wire   [15:0] data_reg;
  tri   [15:0] databus;
  tri   [14:0] addr_out;
  tri   re_out;
  tri   we_out;
  assign databus_out[15] = databus[15];
  assign databus_out[14] = databus[14];
  assign databus_out[13] = databus[13];
  assign databus_out[12] = databus[12];
  assign databus_out[11] = databus[11];
  assign databus_out[10] = databus[10];
  assign databus_out[9] = databus[9];
  assign databus_out[8] = databus[8];
  assign databus_out[7] = databus[7];
  assign databus_out[6] = databus[6];
  assign databus_out[5] = databus[5];
  assign databus_out[4] = databus[4];
  assign databus_out[3] = databus[3];
  assign databus_out[2] = databus[2];
  assign databus_out[1] = databus[1];
  assign databus_out[0] = databus[0];

  DFFSR tem_reg ( .D(strb_in), .CLK(clk), .R(rst_n), .S(1'b1), .Q(tem) );
  DFFSR tem2_reg ( .D(tem), .CLK(clk), .R(rst_n), .S(1'b1), .Q(tem2) );
  DFFSR we_reg ( .D(n274), .CLK(clk), .R(rst_n), .S(1'b1), .Q(we) );
  DFFSR \opcode_reg[15]  ( .D(n125), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        opp[15]) );
  DFFSR \state_reg[3]  ( .D(n331), .CLK(clk), .R(rst_n), .S(1'b1), .Q(state[3]) );
  DFFSR \counter_reg[4]  ( .D(n293), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        counter[4]) );
  DFFSR \state_reg[2]  ( .D(n330), .CLK(clk), .R(rst_n), .S(1'b1), .Q(state[2]) );
  DFFSR \state_reg[0]  ( .D(n328), .CLK(clk), .R(rst_n), .S(1'b1), .Q(state[0]) );
  DFFSR \state_reg[1]  ( .D(n329), .CLK(clk), .R(rst_n), .S(1'b1), .Q(state[1]) );
  DFFPOSX1 \data_reg_reg[0]  ( .D(n103), .CLK(clk), .Q(data_reg[0]) );
  DFFPOSX1 \data_reg_reg[1]  ( .D(n70), .CLK(clk), .Q(data_reg[1]) );
  DFFPOSX1 \data_reg_reg[2]  ( .D(n136), .CLK(clk), .Q(data_reg[2]) );
  DFFPOSX1 \data_reg_reg[3]  ( .D(n66), .CLK(clk), .Q(data_reg[3]) );
  DFFPOSX1 \data_reg_reg[4]  ( .D(n145), .CLK(clk), .Q(data_reg[4]) );
  DFFPOSX1 \data_reg_reg[5]  ( .D(n62), .CLK(clk), .Q(data_reg[5]) );
  DFFPOSX1 \data_reg_reg[6]  ( .D(n148), .CLK(clk), .Q(data_reg[6]) );
  DFFPOSX1 \data_reg_reg[7]  ( .D(n58), .CLK(clk), .Q(data_reg[7]) );
  DFFPOSX1 \data_reg_reg[8]  ( .D(n153), .CLK(clk), .Q(data_reg[8]) );
  DFFPOSX1 \data_reg_reg[9]  ( .D(n57), .CLK(clk), .Q(data_reg[9]) );
  DFFPOSX1 \data_reg_reg[10]  ( .D(n92), .CLK(clk), .Q(data_reg[10]) );
  DFFPOSX1 \data_reg_reg[11]  ( .D(n113), .CLK(clk), .Q(data_reg[11]) );
  DFFPOSX1 \data_reg_reg[12]  ( .D(n76), .CLK(clk), .Q(data_reg[12]) );
  DFFPOSX1 \data_reg_reg[13]  ( .D(n118), .CLK(clk), .Q(data_reg[13]) );
  DFFPOSX1 \data_reg_reg[14]  ( .D(n71), .CLK(clk), .Q(data_reg[14]) );
  DFFPOSX1 \data_reg_reg[15]  ( .D(n121), .CLK(clk), .Q(data_reg[15]) );
  DFFSR \opcode_reg[0]  ( .D(n326), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[0])
         );
  DFFSR \opcode_reg[1]  ( .D(n324), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[1])
         );
  DFFSR \opcode_reg[2]  ( .D(n131), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[2])
         );
  DFFSR \opcode_reg[3]  ( .D(n64), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[3])
         );
  DFFSR \opcode_reg[4]  ( .D(n139), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[4])
         );
  DFFSR \opcode_reg[5]  ( .D(n60), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[5])
         );
  DFFSR \opcode_reg[6]  ( .D(n314), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[6])
         );
  DFFSR \opcode_reg[7]  ( .D(n312), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[7])
         );
  DFFSR \opcode_reg[8]  ( .D(n152), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[8])
         );
  DFFSR \opcode_reg[9]  ( .D(n56), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[9])
         );
  DFFSR \opcode_reg[10]  ( .D(n89), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[10]) );
  DFFSR \opcode_reg[11]  ( .D(n106), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        opp[11]) );
  DFFSR \opcode_reg[12]  ( .D(n72), .CLK(clk), .R(rst_n), .S(1'b1), .Q(opp[12]) );
  DFFSR \opcode_reg[13]  ( .D(n300), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        opp[13]) );
  DFFSR \opcode_reg[14]  ( .D(n298), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        opp[14]) );
  DFFSR \counter_reg[3]  ( .D(n294), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        counter[3]) );
  DFFSR \counter_reg[0]  ( .D(n297), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        counter[0]) );
  DFFSR \counter_reg[1]  ( .D(n296), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        counter[1]) );
  DFFSR \counter_reg[2]  ( .D(n295), .CLK(clk), .R(rst_n), .S(1'b1), .Q(
        counter[2]) );
  DFFSR \addr_reg[15]  ( .D(n276), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[15]) );
  DFFSR \addr_reg[0]  ( .D(n291), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[0])
         );
  DFFSR \addr_reg[1]  ( .D(n290), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[1])
         );
  DFFSR \addr_reg[2]  ( .D(n289), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[2])
         );
  DFFSR \addr_reg[3]  ( .D(n288), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[3])
         );
  DFFSR \addr_reg[4]  ( .D(n287), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[4])
         );
  DFFSR \addr_reg[5]  ( .D(n286), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[5])
         );
  DFFSR \addr_reg[6]  ( .D(n285), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[6])
         );
  DFFSR \addr_reg[7]  ( .D(n284), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[7])
         );
  DFFSR \addr_reg[8]  ( .D(n283), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[8])
         );
  DFFSR \addr_reg[9]  ( .D(n282), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[9])
         );
  DFFSR \addr_reg[10]  ( .D(n281), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[10]) );
  DFFSR \addr_reg[11]  ( .D(n280), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[11]) );
  DFFSR \addr_reg[12]  ( .D(n279), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[12]) );
  DFFSR \addr_reg[13]  ( .D(n278), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[13]) );
  DFFSR \addr_reg[14]  ( .D(n277), .CLK(clk), .R(rst_n), .S(1'b1), .Q(addr[14]) );
  DFFSR re_reg ( .D(nextre), .CLK(clk), .R(rst_n), .S(1'b1), .Q(re) );
  NOR2X1 U4 ( .A(n1), .B(n2), .Y(strb_matrix) );
  NOR2X1 U5 ( .A(n2), .B(n3), .Y(strb_cor) );
  OAI21X1 U6 ( .A(n211), .B(n322), .C(n164), .Y(nextre) );
  NAND2X1 U8 ( .A(n7), .B(n8), .Y(n276) );
  AOI22X1 U9 ( .A(addr[15]), .B(n4), .C(N312), .D(n179), .Y(n8) );
  AOI22X1 U10 ( .A(rast_addr[15]), .B(n201), .C(databus[15]), .D(n212), .Y(n7)
         );
  NAND2X1 U11 ( .A(n13), .B(n14), .Y(n277) );
  AOI22X1 U12 ( .A(n4), .B(addr[14]), .C(N311), .D(n179), .Y(n14) );
  AOI22X1 U13 ( .A(rast_addr[14]), .B(n201), .C(databus[14]), .D(n212), .Y(n13) );
  NAND2X1 U14 ( .A(n15), .B(n16), .Y(n278) );
  AOI22X1 U15 ( .A(n4), .B(addr[13]), .C(N310), .D(n179), .Y(n16) );
  AOI22X1 U16 ( .A(rast_addr[13]), .B(n201), .C(databus[13]), .D(n212), .Y(n15) );
  NAND2X1 U17 ( .A(n17), .B(n18), .Y(n279) );
  AOI22X1 U18 ( .A(n4), .B(addr[12]), .C(N309), .D(n179), .Y(n18) );
  AOI22X1 U19 ( .A(rast_addr[12]), .B(n201), .C(databus[12]), .D(n212), .Y(n17) );
  NAND2X1 U20 ( .A(n19), .B(n20), .Y(n280) );
  AOI22X1 U21 ( .A(n4), .B(addr[11]), .C(N308), .D(n179), .Y(n20) );
  AOI22X1 U22 ( .A(rast_addr[11]), .B(n201), .C(databus[11]), .D(n212), .Y(n19) );
  NAND2X1 U23 ( .A(n21), .B(n22), .Y(n281) );
  AOI22X1 U24 ( .A(n4), .B(addr[10]), .C(N307), .D(n179), .Y(n22) );
  AOI22X1 U25 ( .A(rast_addr[10]), .B(n201), .C(databus[10]), .D(n212), .Y(n21) );
  NAND2X1 U26 ( .A(n23), .B(n24), .Y(n282) );
  AOI22X1 U27 ( .A(n4), .B(addr[9]), .C(N306), .D(n179), .Y(n24) );
  AOI22X1 U28 ( .A(rast_addr[9]), .B(n201), .C(databus[9]), .D(n212), .Y(n23)
         );
  NAND2X1 U29 ( .A(n25), .B(n26), .Y(n283) );
  AOI22X1 U30 ( .A(n4), .B(addr[8]), .C(N305), .D(n179), .Y(n26) );
  AOI22X1 U31 ( .A(rast_addr[8]), .B(n201), .C(databus[8]), .D(n212), .Y(n25)
         );
  NAND2X1 U32 ( .A(n27), .B(n28), .Y(n284) );
  AOI22X1 U33 ( .A(n4), .B(addr[7]), .C(N304), .D(n179), .Y(n28) );
  AOI22X1 U34 ( .A(rast_addr[7]), .B(n201), .C(databus[7]), .D(n212), .Y(n27)
         );
  NAND2X1 U35 ( .A(n29), .B(n30), .Y(n285) );
  AOI22X1 U36 ( .A(n4), .B(addr[6]), .C(N303), .D(n179), .Y(n30) );
  AOI22X1 U37 ( .A(rast_addr[6]), .B(n201), .C(databus[6]), .D(n212), .Y(n29)
         );
  NAND2X1 U38 ( .A(n31), .B(n32), .Y(n286) );
  AOI22X1 U39 ( .A(n4), .B(addr[5]), .C(N302), .D(n179), .Y(n32) );
  AOI22X1 U40 ( .A(rast_addr[5]), .B(n201), .C(databus[5]), .D(n212), .Y(n31)
         );
  NAND2X1 U41 ( .A(n33), .B(n34), .Y(n287) );
  AOI22X1 U42 ( .A(n4), .B(addr[4]), .C(N301), .D(n179), .Y(n34) );
  AOI22X1 U43 ( .A(rast_addr[4]), .B(n201), .C(databus[4]), .D(n212), .Y(n33)
         );
  NAND2X1 U44 ( .A(n35), .B(n36), .Y(n288) );
  AOI22X1 U45 ( .A(n4), .B(addr[3]), .C(N300), .D(n179), .Y(n36) );
  AOI22X1 U46 ( .A(rast_addr[3]), .B(n201), .C(databus[3]), .D(n212), .Y(n35)
         );
  NAND2X1 U47 ( .A(n37), .B(n38), .Y(n289) );
  AOI22X1 U48 ( .A(n4), .B(addr[2]), .C(N299), .D(n179), .Y(n38) );
  AOI22X1 U49 ( .A(rast_addr[2]), .B(n201), .C(databus[2]), .D(n212), .Y(n37)
         );
  NAND2X1 U50 ( .A(n39), .B(n40), .Y(n290) );
  AOI22X1 U51 ( .A(n4), .B(addr[1]), .C(N298), .D(n179), .Y(n40) );
  AOI22X1 U52 ( .A(rast_addr[1]), .B(n201), .C(databus[1]), .D(n212), .Y(n39)
         );
  NAND2X1 U53 ( .A(n41), .B(n42), .Y(n291) );
  AOI22X1 U54 ( .A(n4), .B(addr[0]), .C(N297), .D(n179), .Y(n42) );
  NAND3X1 U56 ( .A(n45), .B(n46), .C(n192), .Y(n44) );
  NAND3X1 U58 ( .A(n49), .B(n213), .C(n51), .Y(n43) );
  AOI22X1 U59 ( .A(rast_addr[0]), .B(n201), .C(databus[0]), .D(n212), .Y(n41)
         );
  AOI22X1 U63 ( .A(databus[15]), .B(n11), .C(n5), .D(data_reg[15]), .Y(n54) );
  OAI21X1 U64 ( .A(n188), .B(n217), .C(n59), .Y(n293) );
  NAND2X1 U65 ( .A(N317), .B(n179), .Y(n59) );
  OAI21X1 U66 ( .A(n188), .B(n299), .C(n61), .Y(n294) );
  NAND2X1 U67 ( .A(N316), .B(n179), .Y(n61) );
  OAI21X1 U68 ( .A(n188), .B(n303), .C(n63), .Y(n295) );
  NAND2X1 U69 ( .A(N315), .B(n179), .Y(n63) );
  OAI21X1 U70 ( .A(n188), .B(n302), .C(n65), .Y(n296) );
  NAND2X1 U71 ( .A(N314), .B(n179), .Y(n65) );
  OAI21X1 U72 ( .A(n188), .B(n301), .C(n67), .Y(n297) );
  NAND2X1 U73 ( .A(n301), .B(n179), .Y(n67) );
  NAND3X1 U75 ( .A(n69), .B(n213), .C(n191), .Y(n68) );
  OAI22X1 U77 ( .A(n9), .B(n292), .C(n73), .D(n10), .Y(n298) );
  AOI22X1 U80 ( .A(databus[14]), .B(n11), .C(n5), .D(data_reg[14]), .Y(n75) );
  OAI22X1 U81 ( .A(n9), .B(n275), .C(n77), .D(n10), .Y(n300) );
  AOI22X1 U84 ( .A(databus[13]), .B(n11), .C(n5), .D(data_reg[13]), .Y(n78) );
  AOI22X1 U86 ( .A(n10), .B(opp[12]), .C(databus[12]), .D(n9), .Y(n79) );
  AOI22X1 U88 ( .A(databus[12]), .B(n11), .C(n5), .D(data_reg[12]), .Y(n80) );
  AOI22X1 U90 ( .A(n74), .B(opp[11]), .C(databus[11]), .D(n9), .Y(n81) );
  AOI22X1 U92 ( .A(databus[11]), .B(n11), .C(n5), .D(data_reg[11]), .Y(n82) );
  AOI22X1 U94 ( .A(n74), .B(opp[10]), .C(databus[10]), .D(n9), .Y(n83) );
  AOI22X1 U96 ( .A(databus[10]), .B(n11), .C(n5), .D(data_reg[10]), .Y(n84) );
  AOI22X1 U98 ( .A(n74), .B(opp[9]), .C(databus[9]), .D(n9), .Y(n85) );
  AOI22X1 U100 ( .A(databus[9]), .B(n11), .C(n5), .D(data_reg[9]), .Y(n86) );
  AOI22X1 U102 ( .A(n74), .B(opp[8]), .C(databus[8]), .D(n9), .Y(n87) );
  AOI22X1 U104 ( .A(databus[8]), .B(n11), .C(n5), .D(data_reg[8]), .Y(n88) );
  OAI22X1 U105 ( .A(n9), .B(n227), .C(n90), .D(n10), .Y(n312) );
  AOI22X1 U108 ( .A(databus[7]), .B(n11), .C(n5), .D(data_reg[7]), .Y(n91) );
  OAI22X1 U109 ( .A(n9), .B(n226), .C(n93), .D(n10), .Y(n314) );
  AOI22X1 U112 ( .A(databus[6]), .B(n11), .C(n5), .D(data_reg[6]), .Y(n94) );
  AOI22X1 U114 ( .A(n74), .B(opp[5]), .C(databus[5]), .D(n9), .Y(n95) );
  AOI22X1 U116 ( .A(databus[5]), .B(n11), .C(n5), .D(data_reg[5]), .Y(n96) );
  AOI22X1 U118 ( .A(n74), .B(opp[4]), .C(databus[4]), .D(n9), .Y(n97) );
  AOI22X1 U120 ( .A(databus[4]), .B(n11), .C(n5), .D(data_reg[4]), .Y(n98) );
  AOI22X1 U122 ( .A(n74), .B(opp[3]), .C(databus[3]), .D(n9), .Y(n99) );
  AOI22X1 U124 ( .A(databus[3]), .B(n11), .C(n5), .D(data_reg[3]), .Y(n100) );
  AOI22X1 U126 ( .A(n74), .B(opp[2]), .C(databus[2]), .D(n9), .Y(n101) );
  AOI22X1 U128 ( .A(databus[2]), .B(n11), .C(n5), .D(data_reg[2]), .Y(n102) );
  OAI22X1 U129 ( .A(n9), .B(n224), .C(n104), .D(n10), .Y(n324) );
  AOI22X1 U132 ( .A(databus[1]), .B(n11), .C(n5), .D(data_reg[1]), .Y(n105) );
  OAI22X1 U133 ( .A(n9), .B(n223), .C(n107), .D(n10), .Y(n326) );
  AOI22X1 U136 ( .A(databus[0]), .B(n11), .C(n5), .D(data_reg[0]), .Y(n108) );
  NAND3X1 U139 ( .A(n191), .B(n69), .C(rst_n), .Y(n110) );
  NAND3X1 U140 ( .A(n46), .B(n2), .C(n111), .Y(n109) );
  OAI21X1 U141 ( .A(n112), .B(n221), .C(n114), .Y(n328) );
  OAI21X1 U142 ( .A(n115), .B(n116), .C(n112), .Y(n114) );
  OAI21X1 U143 ( .A(n117), .B(n46), .C(n181), .Y(n116) );
  NAND2X1 U145 ( .A(n120), .B(n111), .Y(n115) );
  OAI21X1 U146 ( .A(n112), .B(n222), .C(n122), .Y(n329) );
  OAI21X1 U147 ( .A(n123), .B(n124), .C(n112), .Y(n122) );
  NAND2X1 U148 ( .A(n45), .B(n211), .Y(n124) );
  NOR2X1 U149 ( .A(n216), .B(n126), .Y(n45) );
  OAI21X1 U150 ( .A(n127), .B(n128), .C(n129), .Y(n126) );
  NAND2X1 U152 ( .A(n130), .B(n218), .Y(n69) );
  NAND3X1 U153 ( .A(n132), .B(n133), .C(n134), .Y(n330) );
  NOR2X1 U154 ( .A(n123), .B(n135), .Y(n134) );
  OAI21X1 U155 ( .A(n112), .B(n220), .C(n120), .Y(n135) );
  NAND3X1 U157 ( .A(counter[2]), .B(counter[1]), .C(n215), .Y(n138) );
  NAND3X1 U159 ( .A(n299), .B(n217), .C(n140), .Y(n137) );
  NOR2X1 U160 ( .A(counter[0]), .B(n3), .Y(n140) );
  OAI21X1 U162 ( .A(err), .B(n141), .C(n142), .Y(n123) );
  AOI21X1 U164 ( .A(n144), .B(n164), .C(n12), .Y(n331) );
  NOR2X1 U166 ( .A(n146), .B(n147), .Y(n112) );
  OAI22X1 U167 ( .A(n211), .B(rast_strb), .C(n129), .D(n47), .Y(n147) );
  OAI22X1 U169 ( .A(n133), .B(n333), .C(n141), .D(math_done), .Y(n146) );
  OAI21X1 U171 ( .A(n49), .B(n151), .C(n51), .Y(n150) );
  OAI21X1 U172 ( .A(n168), .B(n175), .C(n154), .Y(n151) );
  NAND3X1 U173 ( .A(n301), .B(n299), .C(n155), .Y(n154) );
  OAI21X1 U174 ( .A(n156), .B(n157), .C(n158), .Y(n155) );
  NAND3X1 U175 ( .A(counter[2]), .B(counter[1]), .C(n159), .Y(n158) );
  NOR2X1 U176 ( .A(counter[4]), .B(n3), .Y(n159) );
  NAND2X1 U177 ( .A(counter[4]), .B(n175), .Y(n157) );
  NAND2X1 U178 ( .A(n302), .B(n303), .Y(n156) );
  NAND3X1 U184 ( .A(n160), .B(n224), .C(opp[0]), .Y(n1) );
  NAND3X1 U187 ( .A(n160), .B(n223), .C(opp[1]), .Y(n3) );
  NOR2X1 U190 ( .A(n163), .B(n225), .Y(n162) );
  NOR3X1 U192 ( .A(opp[4]), .B(opp[5]), .C(opp[3]), .Y(n165) );
  NAND3X1 U193 ( .A(n226), .B(n227), .C(n166), .Y(n163) );
  NOR2X1 U194 ( .A(opp[9]), .B(opp[8]), .Y(n166) );
  NOR2X1 U197 ( .A(n167), .B(n228), .Y(n161) );
  NOR3X1 U199 ( .A(opp[11]), .B(opp[12]), .C(opp[10]), .Y(n169) );
  NAND3X1 U200 ( .A(n275), .B(n292), .C(n170), .Y(n167) );
  NOR2X1 U201 ( .A(opp[2]), .B(opp[15]), .Y(n170) );
  NOR2X1 U204 ( .A(n274), .B(n149), .Y(n144) );
  NOR2X1 U205 ( .A(rast_done), .B(n53), .Y(n149) );
  AOI22X1 U207 ( .A(n10), .B(opp[15]), .C(databus[15]), .D(n9), .Y(n171) );
  NAND3X1 U209 ( .A(n191), .B(n46), .C(n132), .Y(n74) );
  NOR2X1 U210 ( .A(n274), .B(n179), .Y(n132) );
  NAND3X1 U212 ( .A(n218), .B(n222), .C(state[3]), .Y(n2) );
  NAND3X1 U214 ( .A(n53), .B(n49), .C(n173), .Y(n172) );
  NOR2X1 U215 ( .A(n48), .B(n119), .Y(n173) );
  NAND3X1 U216 ( .A(n52), .B(n51), .C(n129), .Y(n119) );
  NAND2X1 U217 ( .A(n174), .B(n219), .Y(n129) );
  NAND2X1 U218 ( .A(n219), .B(state[3]), .Y(n51) );
  NAND2X1 U219 ( .A(n174), .B(n218), .Y(n52) );
  NAND3X1 U221 ( .A(n141), .B(n143), .C(n133), .Y(n48) );
  NAND3X1 U222 ( .A(state[2]), .B(state[0]), .C(n174), .Y(n133) );
  NAND3X1 U223 ( .A(state[3]), .B(n177), .C(state[2]), .Y(n143) );
  XOR2X1 U224 ( .A(state[1]), .B(state[0]), .Y(n177) );
  NAND3X1 U225 ( .A(n130), .B(n221), .C(state[2]), .Y(n49) );
  NAND3X1 U226 ( .A(state[2]), .B(n221), .C(n174), .Y(n53) );
  NOR2X1 U227 ( .A(n222), .B(state[3]), .Y(n174) );
  OAI21X1 U229 ( .A(n176), .B(n128), .C(n111), .Y(n274) );
  NAND3X1 U230 ( .A(state[2]), .B(state[3]), .C(n178), .Y(n111) );
  NOR2X1 U231 ( .A(state[1]), .B(state[0]), .Y(n178) );
  NAND2X1 U232 ( .A(state[1]), .B(state[3]), .Y(n128) );
  NAND2X1 U233 ( .A(state[0]), .B(n220), .Y(n176) );
  NOR2X1 U235 ( .A(n332), .B(n180), .Y(init_rast) );
  NAND3X1 U237 ( .A(n130), .B(state[0]), .C(state[2]), .Y(n141) );
  NOR2X1 U239 ( .A(n47), .B(n46), .Y(gpu_done) );
  NAND2X1 U240 ( .A(n130), .B(n219), .Y(n46) );
  NAND2X1 U242 ( .A(n220), .B(n221), .Y(n127) );
  NOR2X1 U245 ( .A(state[3]), .B(state[1]), .Y(n130) );
  NAND2X1 U247 ( .A(tem), .B(n50), .Y(n117) );
  AOI21X1 U249 ( .A(n182), .B(n183), .C(data_reg[9]), .Y(n200) );
  AOI21X1 U250 ( .A(n184), .B(n182), .C(data_reg[8]), .Y(n202) );
  AOI21X1 U251 ( .A(n185), .B(n186), .C(data_reg[7]), .Y(n203) );
  AOI21X1 U252 ( .A(n187), .B(n186), .C(data_reg[6]), .Y(n204) );
  AOI21X1 U253 ( .A(n186), .B(n183), .C(data_reg[5]), .Y(n205) );
  AOI21X1 U254 ( .A(n186), .B(n184), .C(data_reg[4]), .Y(n206) );
  NOR2X1 U255 ( .A(n323), .B(rast_index[3]), .Y(n186) );
  AOI21X1 U256 ( .A(n189), .B(n185), .C(data_reg[3]), .Y(n207) );
  AOI21X1 U257 ( .A(n189), .B(n187), .C(data_reg[2]), .Y(n208) );
  AOI21X1 U258 ( .A(n189), .B(n183), .C(data_reg[1]), .Y(n209) );
  AOI21X1 U259 ( .A(n190), .B(n185), .C(data_reg[15]), .Y(n194) );
  AOI21X1 U260 ( .A(n190), .B(n187), .C(data_reg[14]), .Y(n195) );
  AOI21X1 U261 ( .A(n190), .B(n183), .C(data_reg[13]), .Y(n196) );
  NOR2X1 U262 ( .A(n327), .B(rast_index[1]), .Y(n183) );
  AOI21X1 U263 ( .A(n190), .B(n184), .C(data_reg[12]), .Y(n197) );
  NOR2X1 U264 ( .A(n323), .B(n325), .Y(n190) );
  AOI21X1 U266 ( .A(n185), .B(n182), .C(data_reg[11]), .Y(n198) );
  AOI21X1 U268 ( .A(n187), .B(n182), .C(data_reg[10]), .Y(n199) );
  NOR2X1 U269 ( .A(n325), .B(rast_index[2]), .Y(n182) );
  NAND3X1 U274 ( .A(n333), .B(n321), .C(we), .Y(n193) );
  AOI21X1 U276 ( .A(n189), .B(n184), .C(data_reg[0]), .Y(n210) );
  NOR2X1 U277 ( .A(rast_index[1]), .B(rast_index[0]), .Y(n184) );
  NOR2X1 U278 ( .A(rast_index[3]), .B(rast_index[2]), .Y(n189) );
  INVX2 U78 ( .A(databus[14]), .Y(n73) );
  INVX2 U82 ( .A(databus[13]), .Y(n77) );
  INVX2 U106 ( .A(databus[7]), .Y(n90) );
  INVX2 U110 ( .A(databus[6]), .Y(n93) );
  INVX2 U130 ( .A(databus[1]), .Y(n104) );
  INVX2 U134 ( .A(databus[0]), .Y(n107) );
  OR2X2 U156 ( .A(n137), .B(n138), .Y(n120) );
  AND2X2 U163 ( .A(n143), .B(n52), .Y(n142) );
  AND2X2 U189 ( .A(n161), .B(n162), .Y(n160) );
  OR2X2 U236 ( .A(n141), .B(err), .Y(n180) );
  AND2X2 U267 ( .A(rast_index[1]), .B(rast_index[0]), .Y(n185) );
  AND2X2 U271 ( .A(rast_index[1]), .B(n327), .Y(n187) );
  gpu_controller_DW01_inc_1 add_212 ( .A(addr), .SUM({N312, N311, N310, N309, 
        N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297}) );
  HAX1 \add_213/U1_1_1  ( .A(counter[1]), .B(counter[0]), .YC(
        \add_213/carry[2] ), .YS(N314) );
  HAX1 \add_213/U1_1_2  ( .A(counter[2]), .B(\add_213/carry[2] ), .YC(
        \add_213/carry[3] ), .YS(N315) );
  HAX1 \add_213/U1_1_3  ( .A(counter[3]), .B(\add_213/carry[3] ), .YC(
        \add_213/carry[4] ), .YS(N316) );
  TBUFX1 \databus_tri[15]  ( .A(n194), .EN(n6), .Y(databus[15]) );
  TBUFX1 \databus_tri[14]  ( .A(n195), .EN(n6), .Y(databus[14]) );
  TBUFX1 \databus_tri[2]  ( .A(n208), .EN(n6), .Y(databus[2]) );
  TBUFX1 \databus_tri[3]  ( .A(n207), .EN(n6), .Y(databus[3]) );
  TBUFX1 \databus_tri[4]  ( .A(n206), .EN(n6), .Y(databus[4]) );
  TBUFX1 \databus_tri[12]  ( .A(n197), .EN(n6), .Y(databus[12]) );
  TBUFX1 \databus_tri[8]  ( .A(n202), .EN(n6), .Y(databus[8]) );
  TBUFX1 \databus_tri[10]  ( .A(n199), .EN(n6), .Y(databus[10]) );
  TBUFX1 \databus_tri[11]  ( .A(n198), .EN(n6), .Y(databus[11]) );
  TBUFX1 \databus_tri[0]  ( .A(n210), .EN(n6), .Y(databus[0]) );
  TBUFX1 \databus_tri[5]  ( .A(n205), .EN(n6), .Y(databus[5]) );
  TBUFX1 \databus_tri[9]  ( .A(n200), .EN(n6), .Y(databus[9]) );
  TBUFX1 \databus_tri[6]  ( .A(n204), .EN(n6), .Y(databus[6]) );
  TBUFX1 \databus_tri[7]  ( .A(n203), .EN(n6), .Y(databus[7]) );
  TBUFX1 \databus_tri[1]  ( .A(n209), .EN(n6), .Y(databus[1]) );
  TBUFX1 \databus_tri[13]  ( .A(n196), .EN(n6), .Y(databus[13]) );
  TBUFX1 re_out_tri ( .A(n321), .EN(n333), .Y(re_out) );
  TBUFX1 we_out_tri ( .A(n55), .EN(n333), .Y(we_out) );
  TBUFX1 \addr_out_tri[1]  ( .A(n305), .EN(n333), .Y(addr_out[1]) );
  TBUFX1 \addr_out_tri[2]  ( .A(n306), .EN(n333), .Y(addr_out[2]) );
  TBUFX1 \addr_out_tri[3]  ( .A(n307), .EN(n333), .Y(addr_out[3]) );
  TBUFX1 \addr_out_tri[4]  ( .A(n308), .EN(n333), .Y(addr_out[4]) );
  TBUFX1 \addr_out_tri[5]  ( .A(n309), .EN(n333), .Y(addr_out[5]) );
  TBUFX1 \addr_out_tri[6]  ( .A(n310), .EN(n333), .Y(addr_out[6]) );
  TBUFX1 \addr_out_tri[7]  ( .A(n311), .EN(n333), .Y(addr_out[7]) );
  TBUFX1 \addr_out_tri[8]  ( .A(n313), .EN(n333), .Y(addr_out[8]) );
  TBUFX1 \addr_out_tri[9]  ( .A(n315), .EN(n333), .Y(addr_out[9]) );
  TBUFX1 \addr_out_tri[10]  ( .A(n316), .EN(n333), .Y(addr_out[10]) );
  TBUFX1 \addr_out_tri[11]  ( .A(n317), .EN(n333), .Y(addr_out[11]) );
  TBUFX1 \addr_out_tri[12]  ( .A(n318), .EN(n333), .Y(addr_out[12]) );
  TBUFX1 \addr_out_tri[13]  ( .A(n319), .EN(n333), .Y(addr_out[13]) );
  TBUFX1 \addr_out_tri[14]  ( .A(n320), .EN(n333), .Y(addr_out[14]) );
  TBUFX1 \addr_out_tri[0]  ( .A(n304), .EN(n333), .Y(addr_out[0]) );
  OR2X2 U3 ( .A(n43), .B(n44), .Y(n4) );
  INVX2 U7 ( .A(n9), .Y(n10) );
  INVX2 U55 ( .A(n74), .Y(n9) );
  INVX2 U57 ( .A(n5), .Y(n11) );
  INVX2 U60 ( .A(n52), .Y(n212) );
  INVX2 U61 ( .A(n2), .Y(n179) );
  OR2X2 U62 ( .A(n109), .B(n110), .Y(n5) );
  INVX2 U74 ( .A(n53), .Y(n201) );
  INVX2 U76 ( .A(n193), .Y(n6) );
  INVX2 U79 ( .A(ram_in_use), .Y(n333) );
  XOR2X1 U83 ( .A(\add_213/carry[4] ), .B(counter[4]), .Y(N317) );
  INVX2 U85 ( .A(n112), .Y(n12) );
  INVX2 U87 ( .A(n117), .Y(n47) );
  INVX2 U89 ( .A(tem2), .Y(n50) );
  INVX2 U91 ( .A(we), .Y(n55) );
  INVX2 U93 ( .A(n85), .Y(n56) );
  INVX2 U95 ( .A(n86), .Y(n57) );
  INVX2 U97 ( .A(n91), .Y(n58) );
  INVX2 U99 ( .A(n95), .Y(n60) );
  INVX2 U101 ( .A(n96), .Y(n62) );
  INVX2 U103 ( .A(n99), .Y(n64) );
  INVX2 U107 ( .A(n100), .Y(n66) );
  INVX2 U111 ( .A(n105), .Y(n70) );
  INVX2 U113 ( .A(n75), .Y(n71) );
  INVX2 U115 ( .A(n79), .Y(n72) );
  INVX2 U117 ( .A(n80), .Y(n76) );
  INVX2 U119 ( .A(n83), .Y(n89) );
  INVX2 U121 ( .A(n84), .Y(n92) );
  INVX2 U123 ( .A(n108), .Y(n103) );
  INVX2 U125 ( .A(n81), .Y(n106) );
  INVX2 U127 ( .A(n82), .Y(n113) );
  INVX2 U131 ( .A(n78), .Y(n118) );
  INVX2 U135 ( .A(n54), .Y(n121) );
  INVX2 U137 ( .A(n171), .Y(n125) );
  INVX2 U138 ( .A(n101), .Y(n131) );
  INVX2 U144 ( .A(n102), .Y(n136) );
  INVX2 U151 ( .A(n97), .Y(n139) );
  INVX2 U158 ( .A(n98), .Y(n145) );
  INVX2 U161 ( .A(n94), .Y(n148) );
  INVX2 U165 ( .A(n87), .Y(n152) );
  INVX2 U168 ( .A(n88), .Y(n153) );
  INVX2 U170 ( .A(n150), .Y(n164) );
  INVX2 U179 ( .A(n3), .Y(n168) );
  INVX2 U180 ( .A(n1), .Y(n175) );
  INVX2 U181 ( .A(n119), .Y(n181) );
  INVX2 U182 ( .A(n68), .Y(n188) );
  INVX2 U183 ( .A(n172), .Y(n191) );
  INVX2 U185 ( .A(n48), .Y(n192) );
  INVX2 U186 ( .A(n149), .Y(n211) );
  INVX2 U188 ( .A(n274), .Y(n213) );
  INVX2 U191 ( .A(n141), .Y(init_math) );
  INVX2 U195 ( .A(n49), .Y(n215) );
  INVX2 U196 ( .A(n69), .Y(n216) );
  INVX2 U198 ( .A(counter[4]), .Y(n217) );
  INVX2 U202 ( .A(n176), .Y(n218) );
  INVX2 U203 ( .A(n127), .Y(n219) );
  INVX2 U206 ( .A(state[2]), .Y(n220) );
  INVX2 U208 ( .A(state[0]), .Y(n221) );
  INVX2 U211 ( .A(state[1]), .Y(n222) );
  INVX2 U213 ( .A(opp[0]), .Y(n223) );
  INVX2 U220 ( .A(opp[1]), .Y(n224) );
  INVX2 U228 ( .A(n165), .Y(n225) );
  INVX2 U234 ( .A(opp[6]), .Y(n226) );
  INVX2 U238 ( .A(opp[7]), .Y(n227) );
  INVX2 U241 ( .A(n169), .Y(n228) );
  INVX2 U243 ( .A(opp[13]), .Y(n275) );
  INVX2 U244 ( .A(opp[14]), .Y(n292) );
  INVX2 U246 ( .A(counter[3]), .Y(n299) );
  INVX2 U248 ( .A(counter[0]), .Y(n301) );
  INVX2 U265 ( .A(counter[1]), .Y(n302) );
  INVX2 U270 ( .A(counter[2]), .Y(n303) );
  INVX2 U272 ( .A(addr[0]), .Y(n304) );
  INVX2 U273 ( .A(addr[1]), .Y(n305) );
  INVX2 U275 ( .A(addr[2]), .Y(n306) );
  INVX2 U279 ( .A(addr[3]), .Y(n307) );
  INVX2 U280 ( .A(addr[4]), .Y(n308) );
  INVX2 U281 ( .A(addr[5]), .Y(n309) );
  INVX2 U282 ( .A(addr[6]), .Y(n310) );
  INVX2 U283 ( .A(addr[7]), .Y(n311) );
  INVX2 U284 ( .A(addr[8]), .Y(n313) );
  INVX2 U285 ( .A(addr[9]), .Y(n315) );
  INVX2 U286 ( .A(addr[10]), .Y(n316) );
  INVX2 U287 ( .A(addr[11]), .Y(n317) );
  INVX2 U288 ( .A(addr[12]), .Y(n318) );
  INVX2 U289 ( .A(addr[13]), .Y(n319) );
  INVX2 U290 ( .A(addr[14]), .Y(n320) );
  INVX2 U291 ( .A(re), .Y(n321) );
  INVX2 U292 ( .A(rast_strb), .Y(n322) );
  INVX2 U293 ( .A(rast_index[2]), .Y(n323) );
  INVX2 U294 ( .A(rast_index[3]), .Y(n325) );
  INVX2 U340 ( .A(rast_index[0]), .Y(n327) );
  INVX2 U341 ( .A(math_done), .Y(n332) );
endmodule


module overall ( databus, addr_out, re_out, we_out, strb_in, ram_in_use, 
        gpu_done, clk, rst_n );
  inout [15:0] databus;
  output [14:0] addr_out;
  input strb_in, ram_in_use, clk, rst_n;
  output re_out, we_out, gpu_done;
  wire   math_done, init_math, strb_screen, sel, init_rast, rast_done,
         rast_strb, strb_matrix, strb_cor;
  wire   [47:0] point;
  wire   [63:0] row;
  wire   [7:0] screen_cor;
  wire   [1:0] row_sel;
  wire   [7:0] X0;
  wire   [7:0] X1;
  wire   [7:0] Y0;
  wire   [7:0] Y1;
  wire   [3:0] rast_index;
  wire   [15:0] rast_addr;
  tri   [15:0] databus;
  tri   [14:0] addr_out;
  tri   re_out;
  tri   we_out;
  tri   [15:0] databus_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4;

  matrix_math DUT5 ( .screen_cor(screen_cor), .init_matrix(init_math), .clk(
        clk), .rst_n(rst_n), .row_sel({SYNOPSYS_UNCONNECTED__0, row_sel[0]}), 
        .sel(sel), .math_done(math_done), .strb_screen(strb_screen), .point(
        point), .row(row) );
  Rasterizer DUT4 ( .clk(clk), .X0(X0), .X1(X1), .Y0(Y0), .Y1(Y1), .init_rast(
        init_rast), .RST_N(rst_n), .rast_done(rast_done), .rast_strb(rast_strb), .rast_index(rast_index), .rast_addr({SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, rast_addr[11:0]}) );
  screen_buffer DUT3 ( .clk(clk), .strb_screen(strb_screen), .screen_cor(
        screen_cor), .X0(X0), .X1(X1), .Y0(Y0), .Y1(Y1) );
  world_matrix_buffer DUT2 ( .strb_matrix(strb_matrix), .databus_out(
        databus_out), .clk(clk), .row_sel({1'b0, row_sel[0]}), .row(row) );
  coordinate_buffer DUT1 ( .strb_cor(strb_cor), .databus_out(databus_out), 
        .clk(clk), .sel(sel), .point(point) );
  gpu_controller DUT ( .databus(databus), .strb_in(strb_in), .clk(clk), 
        .rst_n(rst_n), .gpu_done(gpu_done), .ram_in_use(ram_in_use), 
        .rast_done(rast_done), .init_rast(init_rast), .rast_addr({1'b0, 1'b0, 
        1'b0, 1'b0, rast_addr[11:0]}), .rast_strb(rast_strb), .rast_index(
        rast_index), .math_done(math_done), .init_math(init_math), 
        .strb_matrix(strb_matrix), .strb_cor(strb_cor), .err(1'b0), .addr_out(
        addr_out), .re_out(re_out), .we_out(we_out), .databus_out(databus_out)
         );
endmodule

